
//
// Verific Verilog Description of module WES207_top
//

module WES207_top (pll_clk, reset_n, tx_slowclk, led0, led1, SCLK, 
            SSB, MOSI, MISO, gpo_pins, lvds_tx_inst1_DATA);
    input pll_clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input reset_n /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input tx_slowclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output led0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output led1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input SCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input SSB /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MOSI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output MISO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]gpo_pins /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]lvds_tx_inst1_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    
    wire \reg_addr[3] , \reg_addr[2] , \spi_slave_inst/bitcnt[2] , \spi_slave_inst/bitcnt[1] , 
        \spi_slave_inst/sync_tx_en[1] , \reg_addr[1] , \spi_slave_inst/bitcnt[0] , 
        \spi_slave_inst/sync_mosi[1] , n18, n19, rw_out, \reg_addr[0] , 
        \spi_slave_inst/d_o[0] , \rx_d[0] , addr_dv, rxdv, \spi_slave_inst/sync_sclk[0] , 
        \spi_slave_inst/bitcnt[4] , \spi_slave_inst/bitcnt[3] , \spi_slave_inst/sync_ss[0] , 
        \spi_slave_inst/d_o[1] , \spi_slave_inst/d_o[2] , \spi_slave_inst/d_o[3] , 
        \spi_slave_inst/d_o[4] , \spi_slave_inst/d_o[5] , \spi_slave_inst/d_o[6] , 
        \spi_slave_inst/d_o[7] , \rx_d[1] , \rx_d[2] , \rx_d[3] , \rx_d[4] , 
        \rx_d[5] , \rx_d[6] , \rx_d[7] , \spi_slave_inst/sync_sclk[1] , 
        \spi_slave_inst/sync_sclk[2] , \spi_slave_inst/sync_ss[1] , \spi_slave_inst/sync_ss[2] , 
        \data_from_led[7] , \data_from_led[6] , \data_from_led[5] , \data_from_led[4] , 
        \data_from_led[3] , \data_from_led[0] , \data_from_led[2] , \data_from_led[1] , 
        \led_inst/counter[0] , \led_inst/ctr_cfg_reg[0] , \led_inst/counter[1] , 
        \led_inst/counter[2] , \led_inst/counter[3] , \led_inst/counter[4] , 
        \led_inst/counter[5] , \led_inst/counter[6] , \led_inst/counter[7] , 
        \led_inst/counter[8] , \led_inst/counter[9] , \led_inst/counter[10] , 
        \led_inst/counter[11] , \led_inst/counter[12] , \led_inst/counter[13] , 
        \led_inst/counter[14] , \led_inst/counter[15] , \led_inst/counter[16] , 
        \led_inst/counter[17] , \led_inst/counter[18] , \led_inst/counter[19] , 
        \led_inst/counter[20] , \led_inst/counter[21] , \led_inst/counter[22] , 
        \led_inst/counter[23] , \led_inst/ctr_cfg_reg[1] , \led_inst/ctr_cfg_reg[2] , 
        \led_inst/ctr_cfg_reg[3] , \led_inst/ctr_cfg_reg[4] , \led_inst/ctr_cfg_reg[5] , 
        \led_inst/ctr_cfg_reg[6] , \led_inst/ctr_cfg_reg[7] , \i11/fifo_inst/buff[4][5] , 
        \gpo_inst/gp_config_reg[0] , \i11/fifo_inst/buff[4][4] , \gpo_inst/gp_config_reg[1] , 
        \gpo_inst/gp_config_reg[2] , \gpo_inst/gp_config_reg[3] , \gpo_inst/gp_config_reg[4] , 
        \gpo_inst/gp_config_reg[5] , \gpo_inst/gp_config_reg[6] , \gpo_inst/gp_config_reg[7] , 
        \i11/fifo_inst/buff[2][0] , \i11/fifo_inst/buff[2][3] , \i11/fifo_inst/buff[1][7] , 
        \i11/fifo_inst/buff[1][6] , \i11/fifo_inst/buff[1][5] , \i11/fifo_inst/buff[2][2] , 
        \i11/fifo_inst/buff[4][3] , \i11/fifo_inst/buff[2][1] , \i11/fifo_inst/buff[4][2] , 
        \i11/fifo_inst/buff[1][4] , \i11/fifo_inst/buff[4][1] , \i11/fifo_inst/buff[4][0] , 
        \i11/fifo_inst/buff[3][7] , \i11/fifo_inst/buff[3][6] , \i11/fifo_inst/buff[3][5] , 
        \i11/fifo_inst/buff[3][4] , \i11/fifo_inst/buff[3][3] , \i11/fifo_inst/buff[3][2] , 
        \i11/fifo_inst/buff[3][1] , \i11/fifo_inst/buff[3][0] , \i11/fifo_inst/buff[2][7] , 
        \tx_dac_fsm_inst/sym_ctr[0] , \tx_dac_fsm_inst/sym_pos[0] , \tx_dac_fsm_inst/state_reg[0] , 
        n125, \tx_dac_fsm_inst/sym_ctr[1] , \tx_dac_fsm_inst/sym_ctr[2] , 
        \tx_dac_fsm_inst/sym_ctr[3] , \i11/fifo_inst/buff[2][6] , n130, 
        n131, n132, \i11/fifo_inst/buff[2][5] , \tx_dac_fsm_inst/zctr[0] , 
        n135, n136, \tx_dac_fsm_inst/sym_ctr[4] , n138, n139, \tx_dac_fsm_inst/dctr[0] , 
        n141, n142, \tx_dac_fsm_inst/dac_config_reg[0] , \tx_dac_fsm_inst/sym_pos[1] , 
        \tx_dac_fsm_inst/sym_pos[2] , \tx_dac_fsm_inst/sym_pos[3] , \tx_dac_fsm_inst/state_reg[1] , 
        \tx_dac_fsm_inst/state_reg[2] , \tx_dac_fsm_inst/state_reg[3] , 
        n150, n151, n152, n153, \tx_dac_fsm_inst/zctr[1] , \tx_dac_fsm_inst/zctr[2] , 
        \tx_dac_fsm_inst/zctr[3] , \tx_dac_fsm_inst/zctr[4] , \tx_dac_fsm_inst/zctr[5] , 
        \tx_dac_fsm_inst/dctr[1] , \tx_dac_fsm_inst/dctr[2] , \tx_dac_fsm_inst/dctr[3] , 
        \tx_dac_fsm_inst/dctr[4] , \tx_dac_fsm_inst/dctr[5] , \fifo_inst/wr_index[0] , 
        \fifo_inst/rd_index[0] , \fifo_inst/length[0] , \fifo_inst/sync_wr[0] , 
        \fifo_inst/sync_rd[0] , \fifo_inst/buff_head[0] , \fifo_inst/wr_index[1] , 
        \fifo_inst/wr_index[2] , \fifo_inst/wr_index[3] , \fifo_inst/wr_index[4] , 
        \fifo_inst/wr_index[5] , \fifo_inst/wr_index[6] , \fifo_inst/wr_index[7] , 
        \fifo_inst/rd_index[1] , \fifo_inst/rd_index[2] , \fifo_inst/rd_index[3] , 
        \fifo_inst/rd_index[4] , \fifo_inst/rd_index[5] , \fifo_inst/rd_index[6] , 
        \fifo_inst/rd_index[7] , \fifo_inst/length[1] , \fifo_inst/length[2] , 
        \fifo_inst/length[3] , \fifo_inst/length[4] , \fifo_inst/length[5] , 
        \fifo_inst/length[6] , \fifo_inst/length[7] , \fifo_inst/sync_wr[1] , 
        \fifo_inst/sync_rd[1] , \i11/fifo_inst/buff[0][1] , \i11/fifo_inst/buff[0][3] , 
        \i11/fifo_inst/buff[0][5] , \i11/fifo_inst/buff[0][7] , \i11/fifo_inst/buff[1][1] , 
        \i11/fifo_inst/buff[1][3] , \i11/fifo_inst/buff[2][4] , \i11/fifo_inst/buff[0][0] , 
        \i11/fifo_inst/buff[0][2] , \i11/fifo_inst/buff[0][4] , \i11/fifo_inst/buff[0][6] , 
        \i11/fifo_inst/buff[1][0] , \i11/fifo_inst/buff[1][2] , \fifo_inst/buff_head[1] , 
        \fifo_inst/buff_head[2] , \fifo_inst/buff_head[3] , \fifo_inst/buff_head[4] , 
        \fifo_inst/buff_head[5] , \fifo_inst/buff_head[6] , \fifo_inst/buff_head[7] , 
        \i11/fifo_inst/buff[4][6] , \i11/fifo_inst/buff[4][7] , \i11/fifo_inst/buff[5][0] , 
        \i11/fifo_inst/buff[5][1] , \i11/fifo_inst/buff[5][2] , \i11/fifo_inst/buff[5][3] , 
        \i11/fifo_inst/buff[5][4] , \i11/fifo_inst/buff[5][5] , \i11/fifo_inst/buff[5][6] , 
        \i11/fifo_inst/buff[5][7] , \i11/fifo_inst/buff[6][0] , \i11/fifo_inst/buff[6][1] , 
        \i11/fifo_inst/buff[6][2] , \i11/fifo_inst/buff[6][3] , \i11/fifo_inst/buff[6][4] , 
        \i11/fifo_inst/buff[6][5] , \i11/fifo_inst/buff[6][6] , \i11/fifo_inst/buff[6][7] , 
        \i11/fifo_inst/buff[7][0] , \i11/fifo_inst/buff[7][1] , \i11/fifo_inst/buff[7][2] , 
        \i11/fifo_inst/buff[7][3] , \i11/fifo_inst/buff[7][4] , \i11/fifo_inst/buff[7][5] , 
        \i11/fifo_inst/buff[7][6] , \i11/fifo_inst/buff[7][7] , \i11/fifo_inst/buff[8][0] , 
        \i11/fifo_inst/buff[8][1] , \i11/fifo_inst/buff[8][2] , \i11/fifo_inst/buff[8][3] , 
        \i11/fifo_inst/buff[8][4] , \i11/fifo_inst/buff[8][5] , \i11/fifo_inst/buff[8][6] , 
        \i11/fifo_inst/buff[8][7] , \i11/fifo_inst/buff[9][0] , \i11/fifo_inst/buff[9][1] , 
        \i11/fifo_inst/buff[9][2] , \i11/fifo_inst/buff[9][3] , \i11/fifo_inst/buff[9][4] , 
        \i11/fifo_inst/buff[9][5] , \i11/fifo_inst/buff[9][6] , \i11/fifo_inst/buff[9][7] , 
        \i11/fifo_inst/buff[10][0] , \i11/fifo_inst/buff[10][1] , \i11/fifo_inst/buff[10][2] , 
        \i11/fifo_inst/buff[10][3] , \i11/fifo_inst/buff[10][4] , \i11/fifo_inst/buff[10][5] , 
        \i11/fifo_inst/buff[10][6] , \i11/fifo_inst/buff[10][7] , \i11/fifo_inst/buff[11][0] , 
        \i11/fifo_inst/buff[11][1] , \i11/fifo_inst/buff[11][2] , \i11/fifo_inst/buff[11][3] , 
        \i11/fifo_inst/buff[11][4] , \i11/fifo_inst/buff[11][5] , \i11/fifo_inst/buff[11][6] , 
        \i11/fifo_inst/buff[11][7] , \i11/fifo_inst/buff[12][0] , \i11/fifo_inst/buff[12][1] , 
        \i11/fifo_inst/buff[12][2] , \i11/fifo_inst/buff[12][3] , \i11/fifo_inst/buff[12][4] , 
        \i11/fifo_inst/buff[12][5] , \i11/fifo_inst/buff[12][6] , \i11/fifo_inst/buff[12][7] , 
        \i11/fifo_inst/buff[13][0] , \i11/fifo_inst/buff[13][1] , \i11/fifo_inst/buff[13][2] , 
        \i11/fifo_inst/buff[13][3] , \i11/fifo_inst/buff[13][4] , \i11/fifo_inst/buff[13][5] , 
        \i11/fifo_inst/buff[13][6] , \i11/fifo_inst/buff[13][7] , \i11/fifo_inst/buff[14][0] , 
        \i11/fifo_inst/buff[14][1] , \i11/fifo_inst/buff[14][2] , \i11/fifo_inst/buff[14][3] , 
        \i11/fifo_inst/buff[14][4] , \i11/fifo_inst/buff[14][5] , \i11/fifo_inst/buff[14][6] , 
        \i11/fifo_inst/buff[14][7] , \i11/fifo_inst/buff[15][0] , \i11/fifo_inst/buff[15][1] , 
        \i11/fifo_inst/buff[15][2] , \i11/fifo_inst/buff[15][3] , \i11/fifo_inst/buff[15][4] , 
        \i11/fifo_inst/buff[15][5] , \i11/fifo_inst/buff[15][6] , \i11/fifo_inst/buff[15][7] , 
        \i11/fifo_inst/buff[16][0] , \i11/fifo_inst/buff[16][1] , \i11/fifo_inst/buff[16][2] , 
        \i11/fifo_inst/buff[16][3] , \i11/fifo_inst/buff[16][4] , \i11/fifo_inst/buff[16][5] , 
        \i11/fifo_inst/buff[16][6] , \i11/fifo_inst/buff[16][7] , \i11/fifo_inst/buff[17][0] , 
        \i11/fifo_inst/buff[17][1] , \i11/fifo_inst/buff[17][2] , \i11/fifo_inst/buff[17][3] , 
        \i11/fifo_inst/buff[17][4] , \i11/fifo_inst/buff[17][5] , \i11/fifo_inst/buff[17][6] , 
        \i11/fifo_inst/buff[17][7] , \i11/fifo_inst/buff[18][0] , \i11/fifo_inst/buff[18][1] , 
        \i11/fifo_inst/buff[18][2] , \i11/fifo_inst/buff[18][3] , \i11/fifo_inst/buff[18][4] , 
        \i11/fifo_inst/buff[18][5] , \i11/fifo_inst/buff[18][6] , \i11/fifo_inst/buff[18][7] , 
        \i11/fifo_inst/buff[19][0] , \i11/fifo_inst/buff[19][1] , \i11/fifo_inst/buff[19][2] , 
        \i11/fifo_inst/buff[19][3] , \i11/fifo_inst/buff[19][4] , \i11/fifo_inst/buff[19][5] , 
        \i11/fifo_inst/buff[19][6] , \i11/fifo_inst/buff[19][7] , \i11/fifo_inst/buff[20][0] , 
        \i11/fifo_inst/buff[20][1] , \i11/fifo_inst/buff[20][2] , \i11/fifo_inst/buff[20][3] , 
        \i11/fifo_inst/buff[20][4] , \i11/fifo_inst/buff[20][5] , \i11/fifo_inst/buff[20][6] , 
        \i11/fifo_inst/buff[20][7] , \i11/fifo_inst/buff[21][0] , \i11/fifo_inst/buff[21][1] , 
        \i11/fifo_inst/buff[21][2] , \i11/fifo_inst/buff[21][3] , \i11/fifo_inst/buff[21][4] , 
        \i11/fifo_inst/buff[21][5] , \i11/fifo_inst/buff[21][6] , \i11/fifo_inst/buff[21][7] , 
        \i11/fifo_inst/buff[22][0] , \i11/fifo_inst/buff[22][1] , \i11/fifo_inst/buff[22][2] , 
        \i11/fifo_inst/buff[22][3] , \i11/fifo_inst/buff[22][4] , \i11/fifo_inst/buff[22][5] , 
        \i11/fifo_inst/buff[22][6] , \i11/fifo_inst/buff[22][7] , \i11/fifo_inst/buff[23][0] , 
        \i11/fifo_inst/buff[23][1] , \i11/fifo_inst/buff[23][2] , \i11/fifo_inst/buff[23][3] , 
        \i11/fifo_inst/buff[23][4] , \i11/fifo_inst/buff[23][5] , \i11/fifo_inst/buff[23][6] , 
        \i11/fifo_inst/buff[23][7] , \i11/fifo_inst/buff[24][0] , \i11/fifo_inst/buff[24][1] , 
        \i11/fifo_inst/buff[24][2] , \i11/fifo_inst/buff[24][3] , \i11/fifo_inst/buff[24][4] , 
        \i11/fifo_inst/buff[24][5] , \i11/fifo_inst/buff[24][6] , \i11/fifo_inst/buff[24][7] , 
        \i11/fifo_inst/buff[25][0] , \i11/fifo_inst/buff[25][1] , \i11/fifo_inst/buff[25][2] , 
        \i11/fifo_inst/buff[25][3] , \i11/fifo_inst/buff[25][4] , \i11/fifo_inst/buff[25][5] , 
        \i11/fifo_inst/buff[25][6] , \i11/fifo_inst/buff[25][7] , \i11/fifo_inst/buff[26][0] , 
        \i11/fifo_inst/buff[26][1] , \i11/fifo_inst/buff[26][2] , \i11/fifo_inst/buff[26][3] , 
        \i11/fifo_inst/buff[26][4] , \i11/fifo_inst/buff[26][5] , \i11/fifo_inst/buff[26][6] , 
        \i11/fifo_inst/buff[26][7] , \i11/fifo_inst/buff[27][0] , \i11/fifo_inst/buff[27][1] , 
        \i11/fifo_inst/buff[27][2] , \i11/fifo_inst/buff[27][3] , \i11/fifo_inst/buff[27][4] , 
        \i11/fifo_inst/buff[27][5] , \i11/fifo_inst/buff[27][6] , \i11/fifo_inst/buff[27][7] , 
        \i11/fifo_inst/buff[28][0] , \i11/fifo_inst/buff[28][1] , \i11/fifo_inst/buff[28][2] , 
        \i11/fifo_inst/buff[28][3] , \i11/fifo_inst/buff[28][4] , \i11/fifo_inst/buff[28][5] , 
        \i11/fifo_inst/buff[28][6] , \i11/fifo_inst/buff[28][7] , \i11/fifo_inst/buff[29][0] , 
        \i11/fifo_inst/buff[29][1] , \i11/fifo_inst/buff[29][2] , \i11/fifo_inst/buff[29][3] , 
        \i11/fifo_inst/buff[29][4] , \i11/fifo_inst/buff[29][5] , \i11/fifo_inst/buff[29][6] , 
        \i11/fifo_inst/buff[29][7] , \i11/fifo_inst/buff[30][0] , \i11/fifo_inst/buff[30][1] , 
        \i11/fifo_inst/buff[30][2] , \i11/fifo_inst/buff[30][3] , \i11/fifo_inst/buff[30][4] , 
        \i11/fifo_inst/buff[30][5] , \i11/fifo_inst/buff[30][6] , \i11/fifo_inst/buff[30][7] , 
        \i11/fifo_inst/buff[31][0] , \i11/fifo_inst/buff[31][1] , \i11/fifo_inst/buff[31][2] , 
        \i11/fifo_inst/buff[31][3] , \i11/fifo_inst/buff[31][4] , \i11/fifo_inst/buff[31][5] , 
        \i11/fifo_inst/buff[31][6] , \i11/fifo_inst/buff[31][7] , \i11/fifo_inst/buff[32][0] , 
        \i11/fifo_inst/buff[32][1] , \i11/fifo_inst/buff[32][2] , \i11/fifo_inst/buff[32][3] , 
        \i11/fifo_inst/buff[32][4] , \i11/fifo_inst/buff[32][5] , \i11/fifo_inst/buff[32][6] , 
        \i11/fifo_inst/buff[32][7] , \i11/fifo_inst/buff[33][0] , \i11/fifo_inst/buff[33][1] , 
        \i11/fifo_inst/buff[33][2] , \i11/fifo_inst/buff[33][3] , \i11/fifo_inst/buff[33][4] , 
        \i11/fifo_inst/buff[33][5] , \i11/fifo_inst/buff[33][6] , \i11/fifo_inst/buff[33][7] , 
        \i11/fifo_inst/buff[34][0] , \i11/fifo_inst/buff[34][1] , \i11/fifo_inst/buff[34][2] , 
        \i11/fifo_inst/buff[34][3] , \i11/fifo_inst/buff[34][4] , \i11/fifo_inst/buff[34][5] , 
        \i11/fifo_inst/buff[34][6] , \i11/fifo_inst/buff[34][7] , \i11/fifo_inst/buff[35][0] , 
        \i11/fifo_inst/buff[35][1] , \i11/fifo_inst/buff[35][2] , \i11/fifo_inst/buff[35][3] , 
        \i11/fifo_inst/buff[35][4] , \i11/fifo_inst/buff[35][5] , \i11/fifo_inst/buff[35][6] , 
        \i11/fifo_inst/buff[35][7] , \i11/fifo_inst/buff[36][0] , \i11/fifo_inst/buff[36][1] , 
        \i11/fifo_inst/buff[36][2] , \i11/fifo_inst/buff[36][3] , \i11/fifo_inst/buff[36][4] , 
        \i11/fifo_inst/buff[36][5] , \i11/fifo_inst/buff[36][6] , \i11/fifo_inst/buff[36][7] , 
        \i11/fifo_inst/buff[37][0] , \i11/fifo_inst/buff[37][1] , \i11/fifo_inst/buff[37][2] , 
        \i11/fifo_inst/buff[37][3] , \i11/fifo_inst/buff[37][4] , \i11/fifo_inst/buff[37][5] , 
        \i11/fifo_inst/buff[37][6] , \i11/fifo_inst/buff[37][7] , \i11/fifo_inst/buff[38][0] , 
        \i11/fifo_inst/buff[38][1] , \i11/fifo_inst/buff[38][2] , \i11/fifo_inst/buff[38][3] , 
        \i11/fifo_inst/buff[38][4] , \i11/fifo_inst/buff[38][5] , \i11/fifo_inst/buff[38][6] , 
        \i11/fifo_inst/buff[38][7] , \i11/fifo_inst/buff[39][0] , \i11/fifo_inst/buff[39][1] , 
        \i11/fifo_inst/buff[39][2] , \i11/fifo_inst/buff[39][3] , \i11/fifo_inst/buff[39][4] , 
        \i11/fifo_inst/buff[39][5] , \i11/fifo_inst/buff[39][6] , \i11/fifo_inst/buff[39][7] , 
        \i11/fifo_inst/buff[40][0] , \i11/fifo_inst/buff[40][1] , \i11/fifo_inst/buff[40][2] , 
        \i11/fifo_inst/buff[40][3] , \i11/fifo_inst/buff[40][4] , \i11/fifo_inst/buff[40][5] , 
        \i11/fifo_inst/buff[40][6] , \i11/fifo_inst/buff[40][7] , \i11/fifo_inst/buff[41][0] , 
        \i11/fifo_inst/buff[41][1] , \i11/fifo_inst/buff[41][2] , \i11/fifo_inst/buff[41][3] , 
        \i11/fifo_inst/buff[41][4] , \i11/fifo_inst/buff[41][5] , \i11/fifo_inst/buff[41][6] , 
        \i11/fifo_inst/buff[41][7] , \i11/fifo_inst/buff[42][0] , \i11/fifo_inst/buff[42][1] , 
        \i11/fifo_inst/buff[42][2] , \i11/fifo_inst/buff[42][3] , \i11/fifo_inst/buff[42][4] , 
        \i11/fifo_inst/buff[42][5] , \i11/fifo_inst/buff[42][6] , \i11/fifo_inst/buff[42][7] , 
        \i11/fifo_inst/buff[43][0] , \i11/fifo_inst/buff[43][1] , \i11/fifo_inst/buff[43][2] , 
        \i11/fifo_inst/buff[43][3] , \i11/fifo_inst/buff[43][4] , \i11/fifo_inst/buff[43][5] , 
        \i11/fifo_inst/buff[43][6] , \i11/fifo_inst/buff[43][7] , \i11/fifo_inst/buff[44][0] , 
        \i11/fifo_inst/buff[44][1] , \i11/fifo_inst/buff[44][2] , \i11/fifo_inst/buff[44][3] , 
        \i11/fifo_inst/buff[44][4] , \i11/fifo_inst/buff[44][5] , \i11/fifo_inst/buff[44][6] , 
        \i11/fifo_inst/buff[44][7] , \i11/fifo_inst/buff[45][0] , \i11/fifo_inst/buff[45][1] , 
        \i11/fifo_inst/buff[45][2] , \i11/fifo_inst/buff[45][3] , \i11/fifo_inst/buff[45][4] , 
        \i11/fifo_inst/buff[45][5] , \i11/fifo_inst/buff[45][6] , \i11/fifo_inst/buff[45][7] , 
        \i11/fifo_inst/buff[46][0] , \i11/fifo_inst/buff[46][1] , \i11/fifo_inst/buff[46][2] , 
        \i11/fifo_inst/buff[46][3] , \i11/fifo_inst/buff[46][4] , \i11/fifo_inst/buff[46][5] , 
        \i11/fifo_inst/buff[46][6] , \i11/fifo_inst/buff[46][7] , \i11/fifo_inst/buff[47][0] , 
        \i11/fifo_inst/buff[47][1] , \i11/fifo_inst/buff[47][2] , \i11/fifo_inst/buff[47][3] , 
        \i11/fifo_inst/buff[47][4] , \i11/fifo_inst/buff[47][5] , \i11/fifo_inst/buff[47][6] , 
        \i11/fifo_inst/buff[47][7] , \i11/fifo_inst/buff[48][0] , \i11/fifo_inst/buff[48][1] , 
        \i11/fifo_inst/buff[48][2] , \i11/fifo_inst/buff[48][3] , \i11/fifo_inst/buff[48][4] , 
        \i11/fifo_inst/buff[48][5] , \i11/fifo_inst/buff[48][6] , \i11/fifo_inst/buff[48][7] , 
        \i11/fifo_inst/buff[49][0] , \i11/fifo_inst/buff[49][1] , \i11/fifo_inst/buff[49][2] , 
        \i11/fifo_inst/buff[49][3] , \i11/fifo_inst/buff[49][4] , \i11/fifo_inst/buff[49][5] , 
        \i11/fifo_inst/buff[49][6] , \i11/fifo_inst/buff[49][7] , \i11/fifo_inst/buff[50][0] , 
        \i11/fifo_inst/buff[50][1] , \i11/fifo_inst/buff[50][2] , \i11/fifo_inst/buff[50][3] , 
        \i11/fifo_inst/buff[50][4] , \i11/fifo_inst/buff[50][5] , \i11/fifo_inst/buff[50][6] , 
        \i11/fifo_inst/buff[50][7] , \i11/fifo_inst/buff[51][0] , \i11/fifo_inst/buff[51][1] , 
        \i11/fifo_inst/buff[51][2] , \i11/fifo_inst/buff[51][3] , \i11/fifo_inst/buff[51][4] , 
        \i11/fifo_inst/buff[51][5] , \i11/fifo_inst/buff[51][6] , \i11/fifo_inst/buff[51][7] , 
        \i11/fifo_inst/buff[52][0] , \i11/fifo_inst/buff[52][1] , \i11/fifo_inst/buff[52][2] , 
        \i11/fifo_inst/buff[52][3] , \i11/fifo_inst/buff[52][4] , \i11/fifo_inst/buff[52][5] , 
        \i11/fifo_inst/buff[52][6] , \i11/fifo_inst/buff[52][7] , \i11/fifo_inst/buff[53][0] , 
        \i11/fifo_inst/buff[53][1] , \i11/fifo_inst/buff[53][2] , \i11/fifo_inst/buff[53][3] , 
        \i11/fifo_inst/buff[53][4] , \i11/fifo_inst/buff[53][5] , \i11/fifo_inst/buff[53][6] , 
        \i11/fifo_inst/buff[53][7] , \i11/fifo_inst/buff[54][0] , \i11/fifo_inst/buff[54][1] , 
        \i11/fifo_inst/buff[54][2] , \i11/fifo_inst/buff[54][3] , \i11/fifo_inst/buff[54][4] , 
        \i11/fifo_inst/buff[54][5] , \i11/fifo_inst/buff[54][6] , \i11/fifo_inst/buff[54][7] , 
        \i11/fifo_inst/buff[55][0] , \i11/fifo_inst/buff[55][1] , \i11/fifo_inst/buff[55][2] , 
        \i11/fifo_inst/buff[55][3] , \i11/fifo_inst/buff[55][4] , \i11/fifo_inst/buff[55][5] , 
        \i11/fifo_inst/buff[55][6] , \i11/fifo_inst/buff[55][7] , \i11/fifo_inst/buff[56][0] , 
        \i11/fifo_inst/buff[56][1] , \i11/fifo_inst/buff[56][2] , \i11/fifo_inst/buff[56][3] , 
        \i11/fifo_inst/buff[56][4] , \i11/fifo_inst/buff[56][5] , \i11/fifo_inst/buff[56][6] , 
        \i11/fifo_inst/buff[56][7] , \i11/fifo_inst/buff[57][0] , \i11/fifo_inst/buff[57][1] , 
        \i11/fifo_inst/buff[57][2] , \i11/fifo_inst/buff[57][3] , \i11/fifo_inst/buff[57][4] , 
        \i11/fifo_inst/buff[57][5] , \i11/fifo_inst/buff[57][6] , \i11/fifo_inst/buff[57][7] , 
        \i11/fifo_inst/buff[58][0] , \i11/fifo_inst/buff[58][1] , \i11/fifo_inst/buff[58][2] , 
        \i11/fifo_inst/buff[58][3] , \i11/fifo_inst/buff[58][4] , \i11/fifo_inst/buff[58][5] , 
        \i11/fifo_inst/buff[58][6] , \i11/fifo_inst/buff[58][7] , \i11/fifo_inst/buff[59][0] , 
        \i11/fifo_inst/buff[59][1] , \i11/fifo_inst/buff[59][2] , \i11/fifo_inst/buff[59][3] , 
        \i11/fifo_inst/buff[59][4] , \i11/fifo_inst/buff[59][5] , \i11/fifo_inst/buff[59][6] , 
        \i11/fifo_inst/buff[59][7] , \i11/fifo_inst/buff[60][0] , \i11/fifo_inst/buff[60][1] , 
        \i11/fifo_inst/buff[60][2] , \i11/fifo_inst/buff[60][3] , \i11/fifo_inst/buff[60][4] , 
        \i11/fifo_inst/buff[60][5] , \i11/fifo_inst/buff[60][6] , \i11/fifo_inst/buff[60][7] , 
        \i11/fifo_inst/buff[61][0] , \i11/fifo_inst/buff[61][1] , \i11/fifo_inst/buff[61][2] , 
        \i11/fifo_inst/buff[61][3] , \i11/fifo_inst/buff[61][4] , \i11/fifo_inst/buff[61][5] , 
        \i11/fifo_inst/buff[61][6] , \i11/fifo_inst/buff[61][7] , \i11/fifo_inst/buff[62][0] , 
        \i11/fifo_inst/buff[62][1] , \i11/fifo_inst/buff[62][2] , \i11/fifo_inst/buff[62][3] , 
        \i11/fifo_inst/buff[62][4] , \i11/fifo_inst/buff[62][5] , \i11/fifo_inst/buff[62][6] , 
        \i11/fifo_inst/buff[62][7] , \i11/fifo_inst/buff[63][0] , \i11/fifo_inst/buff[63][1] , 
        \i11/fifo_inst/buff[63][2] , \i11/fifo_inst/buff[63][3] , \i11/fifo_inst/buff[63][4] , 
        \i11/fifo_inst/buff[63][5] , \i11/fifo_inst/buff[63][6] , \i11/fifo_inst/buff[63][7] , 
        \i11/fifo_inst/buff[64][0] , \i11/fifo_inst/buff[64][1] , \i11/fifo_inst/buff[64][2] , 
        \i11/fifo_inst/buff[64][3] , \i11/fifo_inst/buff[64][4] , \i11/fifo_inst/buff[64][5] , 
        \i11/fifo_inst/buff[64][6] , \i11/fifo_inst/buff[64][7] , \i11/fifo_inst/buff[65][0] , 
        \i11/fifo_inst/buff[65][1] , \i11/fifo_inst/buff[65][2] , \i11/fifo_inst/buff[65][3] , 
        \i11/fifo_inst/buff[65][4] , \i11/fifo_inst/buff[65][5] , \i11/fifo_inst/buff[65][6] , 
        \i11/fifo_inst/buff[65][7] , \i11/fifo_inst/buff[66][0] , \i11/fifo_inst/buff[66][1] , 
        \i11/fifo_inst/buff[66][2] , \i11/fifo_inst/buff[66][3] , \i11/fifo_inst/buff[66][4] , 
        \i11/fifo_inst/buff[66][5] , \i11/fifo_inst/buff[66][6] , \i11/fifo_inst/buff[66][7] , 
        \i11/fifo_inst/buff[67][0] , \i11/fifo_inst/buff[67][1] , \i11/fifo_inst/buff[67][2] , 
        \i11/fifo_inst/buff[67][3] , \i11/fifo_inst/buff[67][4] , \i11/fifo_inst/buff[67][5] , 
        \i11/fifo_inst/buff[67][6] , \i11/fifo_inst/buff[67][7] , \i11/fifo_inst/buff[68][0] , 
        \i11/fifo_inst/buff[68][1] , \i11/fifo_inst/buff[68][2] , \i11/fifo_inst/buff[68][3] , 
        \i11/fifo_inst/buff[68][4] , \i11/fifo_inst/buff[68][5] , \i11/fifo_inst/buff[68][6] , 
        \i11/fifo_inst/buff[68][7] , \i11/fifo_inst/buff[69][0] , \i11/fifo_inst/buff[69][1] , 
        \i11/fifo_inst/buff[69][2] , \i11/fifo_inst/buff[69][3] , \i11/fifo_inst/buff[69][4] , 
        \i11/fifo_inst/buff[69][5] , \i11/fifo_inst/buff[69][6] , \i11/fifo_inst/buff[69][7] , 
        \i11/fifo_inst/buff[70][0] , \i11/fifo_inst/buff[70][1] , \i11/fifo_inst/buff[70][2] , 
        \i11/fifo_inst/buff[70][3] , \i11/fifo_inst/buff[70][4] , \i11/fifo_inst/buff[70][5] , 
        \i11/fifo_inst/buff[70][6] , \i11/fifo_inst/buff[70][7] , \i11/fifo_inst/buff[71][0] , 
        \i11/fifo_inst/buff[71][1] , \i11/fifo_inst/buff[71][2] , \i11/fifo_inst/buff[71][3] , 
        \i11/fifo_inst/buff[71][4] , \i11/fifo_inst/buff[71][5] , \i11/fifo_inst/buff[71][6] , 
        \i11/fifo_inst/buff[71][7] , \i11/fifo_inst/buff[72][0] , \i11/fifo_inst/buff[72][1] , 
        \i11/fifo_inst/buff[72][2] , \i11/fifo_inst/buff[72][3] , \i11/fifo_inst/buff[72][4] , 
        \i11/fifo_inst/buff[72][5] , \i11/fifo_inst/buff[72][6] , \i11/fifo_inst/buff[72][7] , 
        \i11/fifo_inst/buff[73][0] , \i11/fifo_inst/buff[73][1] , \i11/fifo_inst/buff[73][2] , 
        \i11/fifo_inst/buff[73][3] , \i11/fifo_inst/buff[73][4] , \i11/fifo_inst/buff[73][5] , 
        \i11/fifo_inst/buff[73][6] , \i11/fifo_inst/buff[73][7] , \i11/fifo_inst/buff[74][0] , 
        \i11/fifo_inst/buff[74][1] , \i11/fifo_inst/buff[74][2] , \i11/fifo_inst/buff[74][3] , 
        \i11/fifo_inst/buff[74][4] , \i11/fifo_inst/buff[74][5] , \i11/fifo_inst/buff[74][6] , 
        \i11/fifo_inst/buff[74][7] , \i11/fifo_inst/buff[75][0] , \i11/fifo_inst/buff[75][1] , 
        \i11/fifo_inst/buff[75][2] , \i11/fifo_inst/buff[75][3] , \i11/fifo_inst/buff[75][4] , 
        \i11/fifo_inst/buff[75][5] , \i11/fifo_inst/buff[75][6] , \i11/fifo_inst/buff[75][7] , 
        \i11/fifo_inst/buff[76][0] , \i11/fifo_inst/buff[76][1] , \i11/fifo_inst/buff[76][2] , 
        \i11/fifo_inst/buff[76][3] , \i11/fifo_inst/buff[76][4] , \i11/fifo_inst/buff[76][5] , 
        \i11/fifo_inst/buff[76][6] , \i11/fifo_inst/buff[76][7] , \i11/fifo_inst/buff[77][0] , 
        \i11/fifo_inst/buff[77][1] , \i11/fifo_inst/buff[77][2] , \i11/fifo_inst/buff[77][3] , 
        \i11/fifo_inst/buff[77][4] , \i11/fifo_inst/buff[77][5] , \i11/fifo_inst/buff[77][6] , 
        \i11/fifo_inst/buff[77][7] , \i11/fifo_inst/buff[78][0] , \i11/fifo_inst/buff[78][1] , 
        \i11/fifo_inst/buff[78][2] , \i11/fifo_inst/buff[78][3] , \i11/fifo_inst/buff[78][4] , 
        \i11/fifo_inst/buff[78][5] , \i11/fifo_inst/buff[78][6] , \i11/fifo_inst/buff[78][7] , 
        \i11/fifo_inst/buff[79][0] , \i11/fifo_inst/buff[79][1] , \i11/fifo_inst/buff[79][2] , 
        \i11/fifo_inst/buff[79][3] , \i11/fifo_inst/buff[79][4] , \i11/fifo_inst/buff[79][5] , 
        \i11/fifo_inst/buff[79][6] , \i11/fifo_inst/buff[79][7] , \i11/fifo_inst/buff[80][0] , 
        \i11/fifo_inst/buff[80][1] , \i11/fifo_inst/buff[80][2] , \i11/fifo_inst/buff[80][3] , 
        \i11/fifo_inst/buff[80][4] , \i11/fifo_inst/buff[80][5] , \i11/fifo_inst/buff[80][6] , 
        \i11/fifo_inst/buff[80][7] , \i11/fifo_inst/buff[81][0] , \i11/fifo_inst/buff[81][1] , 
        \i11/fifo_inst/buff[81][2] , \i11/fifo_inst/buff[81][3] , \i11/fifo_inst/buff[81][4] , 
        \i11/fifo_inst/buff[81][5] , \i11/fifo_inst/buff[81][6] , \i11/fifo_inst/buff[81][7] , 
        \i11/fifo_inst/buff[82][0] , \i11/fifo_inst/buff[82][1] , \i11/fifo_inst/buff[82][2] , 
        \i11/fifo_inst/buff[82][3] , \i11/fifo_inst/buff[82][4] , \i11/fifo_inst/buff[82][5] , 
        \i11/fifo_inst/buff[82][6] , \i11/fifo_inst/buff[82][7] , \i11/fifo_inst/buff[83][0] , 
        \i11/fifo_inst/buff[83][1] , \i11/fifo_inst/buff[83][2] , \i11/fifo_inst/buff[83][3] , 
        \i11/fifo_inst/buff[83][4] , \i11/fifo_inst/buff[83][5] , \i11/fifo_inst/buff[83][6] , 
        \i11/fifo_inst/buff[83][7] , \i11/fifo_inst/buff[84][0] , \i11/fifo_inst/buff[84][1] , 
        \i11/fifo_inst/buff[84][2] , \i11/fifo_inst/buff[84][3] , \i11/fifo_inst/buff[84][4] , 
        \i11/fifo_inst/buff[84][5] , \i11/fifo_inst/buff[84][6] , \i11/fifo_inst/buff[84][7] , 
        \i11/fifo_inst/buff[85][0] , \i11/fifo_inst/buff[85][1] , \i11/fifo_inst/buff[85][2] , 
        \i11/fifo_inst/buff[85][3] , \i11/fifo_inst/buff[85][4] , \i11/fifo_inst/buff[85][5] , 
        \i11/fifo_inst/buff[85][6] , \i11/fifo_inst/buff[85][7] , \i11/fifo_inst/buff[86][0] , 
        \i11/fifo_inst/buff[86][1] , \i11/fifo_inst/buff[86][2] , \i11/fifo_inst/buff[86][3] , 
        \i11/fifo_inst/buff[86][4] , \i11/fifo_inst/buff[86][5] , \i11/fifo_inst/buff[86][6] , 
        \i11/fifo_inst/buff[86][7] , \i11/fifo_inst/buff[87][0] , \i11/fifo_inst/buff[87][1] , 
        \i11/fifo_inst/buff[87][2] , \i11/fifo_inst/buff[87][3] , \i11/fifo_inst/buff[87][4] , 
        \i11/fifo_inst/buff[87][5] , \i11/fifo_inst/buff[87][6] , \i11/fifo_inst/buff[87][7] , 
        \i11/fifo_inst/buff[88][0] , \i11/fifo_inst/buff[88][1] , \i11/fifo_inst/buff[88][2] , 
        \i11/fifo_inst/buff[88][3] , \i11/fifo_inst/buff[88][4] , \i11/fifo_inst/buff[88][5] , 
        \i11/fifo_inst/buff[88][6] , \i11/fifo_inst/buff[88][7] , \i11/fifo_inst/buff[89][0] , 
        \i11/fifo_inst/buff[89][1] , \i11/fifo_inst/buff[89][2] , \i11/fifo_inst/buff[89][3] , 
        \i11/fifo_inst/buff[89][4] , \i11/fifo_inst/buff[89][5] , \i11/fifo_inst/buff[89][6] , 
        \i11/fifo_inst/buff[89][7] , \i11/fifo_inst/buff[90][0] , \i11/fifo_inst/buff[90][1] , 
        \i11/fifo_inst/buff[90][2] , \i11/fifo_inst/buff[90][3] , \i11/fifo_inst/buff[90][4] , 
        \i11/fifo_inst/buff[90][5] , \i11/fifo_inst/buff[90][6] , \i11/fifo_inst/buff[90][7] , 
        \i11/fifo_inst/buff[91][0] , \i11/fifo_inst/buff[91][1] , \i11/fifo_inst/buff[91][2] , 
        \i11/fifo_inst/buff[91][3] , \i11/fifo_inst/buff[91][4] , \i11/fifo_inst/buff[91][5] , 
        \i11/fifo_inst/buff[91][6] , \i11/fifo_inst/buff[91][7] , \i11/fifo_inst/buff[92][0] , 
        \i11/fifo_inst/buff[92][1] , \i11/fifo_inst/buff[92][2] , \i11/fifo_inst/buff[92][3] , 
        \i11/fifo_inst/buff[92][4] , \i11/fifo_inst/buff[92][5] , \i11/fifo_inst/buff[92][6] , 
        \i11/fifo_inst/buff[92][7] , \i11/fifo_inst/buff[93][0] , \i11/fifo_inst/buff[93][1] , 
        \i11/fifo_inst/buff[93][2] , \i11/fifo_inst/buff[93][3] , \i11/fifo_inst/buff[93][4] , 
        \i11/fifo_inst/buff[93][5] , \i11/fifo_inst/buff[93][6] , \i11/fifo_inst/buff[93][7] , 
        \i11/fifo_inst/buff[94][0] , \i11/fifo_inst/buff[94][1] , \i11/fifo_inst/buff[94][2] , 
        \i11/fifo_inst/buff[94][3] , \i11/fifo_inst/buff[94][4] , \i11/fifo_inst/buff[94][5] , 
        \i11/fifo_inst/buff[94][6] , \i11/fifo_inst/buff[94][7] , \i11/fifo_inst/buff[95][0] , 
        \i11/fifo_inst/buff[95][1] , \i11/fifo_inst/buff[95][2] , \i11/fifo_inst/buff[95][3] , 
        \i11/fifo_inst/buff[95][4] , \i11/fifo_inst/buff[95][5] , \i11/fifo_inst/buff[95][6] , 
        \i11/fifo_inst/buff[95][7] , \i11/fifo_inst/buff[96][0] , \i11/fifo_inst/buff[96][1] , 
        \i11/fifo_inst/buff[96][2] , \i11/fifo_inst/buff[96][3] , \i11/fifo_inst/buff[96][4] , 
        \i11/fifo_inst/buff[96][5] , \i11/fifo_inst/buff[96][6] , \i11/fifo_inst/buff[96][7] , 
        \i11/fifo_inst/buff[97][0] , \i11/fifo_inst/buff[97][1] , \i11/fifo_inst/buff[97][2] , 
        \i11/fifo_inst/buff[97][3] , \i11/fifo_inst/buff[97][4] , \i11/fifo_inst/buff[97][5] , 
        \i11/fifo_inst/buff[97][6] , \i11/fifo_inst/buff[97][7] , \i11/fifo_inst/buff[98][0] , 
        \i11/fifo_inst/buff[98][1] , \i11/fifo_inst/buff[98][2] , \i11/fifo_inst/buff[98][3] , 
        \i11/fifo_inst/buff[98][4] , \i11/fifo_inst/buff[98][5] , \i11/fifo_inst/buff[98][6] , 
        \i11/fifo_inst/buff[98][7] , \i11/fifo_inst/buff[99][0] , \i11/fifo_inst/buff[99][1] , 
        \i11/fifo_inst/buff[99][2] , \i11/fifo_inst/buff[99][3] , \i11/fifo_inst/buff[99][4] , 
        \i11/fifo_inst/buff[99][5] , \i11/fifo_inst/buff[99][6] , \i11/fifo_inst/buff[99][7] , 
        \i11/fifo_inst/buff[100][0] , \i11/fifo_inst/buff[100][1] , \i11/fifo_inst/buff[100][2] , 
        \i11/fifo_inst/buff[100][3] , \i11/fifo_inst/buff[100][4] , \i11/fifo_inst/buff[100][5] , 
        \i11/fifo_inst/buff[100][6] , \i11/fifo_inst/buff[100][7] , \i11/fifo_inst/buff[101][0] , 
        \i11/fifo_inst/buff[101][1] , \i11/fifo_inst/buff[101][2] , \i11/fifo_inst/buff[101][3] , 
        \i11/fifo_inst/buff[101][4] , \i11/fifo_inst/buff[101][5] , \i11/fifo_inst/buff[101][6] , 
        \i11/fifo_inst/buff[101][7] , \i11/fifo_inst/buff[102][0] , \i11/fifo_inst/buff[102][1] , 
        \i11/fifo_inst/buff[102][2] , \i11/fifo_inst/buff[102][3] , \i11/fifo_inst/buff[102][4] , 
        \i11/fifo_inst/buff[102][5] , \i11/fifo_inst/buff[102][6] , \i11/fifo_inst/buff[102][7] , 
        \i11/fifo_inst/buff[103][0] , \i11/fifo_inst/buff[103][1] , \i11/fifo_inst/buff[103][2] , 
        \i11/fifo_inst/buff[103][3] , \i11/fifo_inst/buff[103][4] , \i11/fifo_inst/buff[103][5] , 
        \i11/fifo_inst/buff[103][6] , \i11/fifo_inst/buff[103][7] , \i11/fifo_inst/buff[104][0] , 
        \i11/fifo_inst/buff[104][1] , \i11/fifo_inst/buff[104][2] , \i11/fifo_inst/buff[104][3] , 
        \i11/fifo_inst/buff[104][4] , \i11/fifo_inst/buff[104][5] , \i11/fifo_inst/buff[104][6] , 
        \i11/fifo_inst/buff[104][7] , \i11/fifo_inst/buff[105][0] , \i11/fifo_inst/buff[105][1] , 
        \i11/fifo_inst/buff[105][2] , \i11/fifo_inst/buff[105][3] , \i11/fifo_inst/buff[105][4] , 
        \i11/fifo_inst/buff[105][5] , \i11/fifo_inst/buff[105][6] , \i11/fifo_inst/buff[105][7] , 
        \i11/fifo_inst/buff[106][0] , \i11/fifo_inst/buff[106][1] , \i11/fifo_inst/buff[106][2] , 
        \i11/fifo_inst/buff[106][3] , \i11/fifo_inst/buff[106][4] , \i11/fifo_inst/buff[106][5] , 
        \i11/fifo_inst/buff[106][6] , \i11/fifo_inst/buff[106][7] , \i11/fifo_inst/buff[107][0] , 
        \i11/fifo_inst/buff[107][1] , \i11/fifo_inst/buff[107][2] , \i11/fifo_inst/buff[107][3] , 
        \i11/fifo_inst/buff[107][4] , \i11/fifo_inst/buff[107][5] , \i11/fifo_inst/buff[107][6] , 
        \i11/fifo_inst/buff[107][7] , \i11/fifo_inst/buff[108][0] , \i11/fifo_inst/buff[108][1] , 
        \i11/fifo_inst/buff[108][2] , \i11/fifo_inst/buff[108][3] , \i11/fifo_inst/buff[108][4] , 
        \i11/fifo_inst/buff[108][5] , \i11/fifo_inst/buff[108][6] , \i11/fifo_inst/buff[108][7] , 
        \i11/fifo_inst/buff[109][0] , \i11/fifo_inst/buff[109][1] , \i11/fifo_inst/buff[109][2] , 
        \i11/fifo_inst/buff[109][3] , \i11/fifo_inst/buff[109][4] , \i11/fifo_inst/buff[109][5] , 
        \i11/fifo_inst/buff[109][6] , \i11/fifo_inst/buff[109][7] , \i11/fifo_inst/buff[110][0] , 
        \i11/fifo_inst/buff[110][1] , \i11/fifo_inst/buff[110][2] , \i11/fifo_inst/buff[110][3] , 
        \i11/fifo_inst/buff[110][4] , \i11/fifo_inst/buff[110][5] , \i11/fifo_inst/buff[110][6] , 
        \i11/fifo_inst/buff[110][7] , \i11/fifo_inst/buff[111][0] , \i11/fifo_inst/buff[111][1] , 
        \i11/fifo_inst/buff[111][2] , \i11/fifo_inst/buff[111][3] , n1067, 
        \i11/fifo_inst/buff[111][4] , \i11/fifo_inst/buff[111][5] , n1070, 
        n1071, \i11/fifo_inst/buff[111][6] , n1073, n1074, \i11/fifo_inst/buff[111][7] , 
        \i11/fifo_inst/buff[112][0] , n1077, n1078, \i11/fifo_inst/buff[112][1] , 
        n1080, n1081, \i11/fifo_inst/buff[112][2] , n1083, n1084, 
        \i11/fifo_inst/buff[112][3] , \i11/fifo_inst/buff[112][4] , \i11/fifo_inst/buff[112][5] , 
        \i11/fifo_inst/buff[112][6] , \i11/fifo_inst/buff[112][7] , n1090, 
        \i11/fifo_inst/buff[113][0] , n1092, n1093, \i11/fifo_inst/buff[113][1] , 
        n1095, n1096, \i11/fifo_inst/buff[113][2] , \i11/fifo_inst/buff[113][3] , 
        \i11/fifo_inst/buff[113][4] , \i11/fifo_inst/buff[113][5] , \i11/fifo_inst/buff[113][6] , 
        \i11/fifo_inst/buff[113][7] , \i11/fifo_inst/buff[114][0] , \i11/fifo_inst/buff[114][1] , 
        \i11/fifo_inst/buff[114][2] , \i11/fifo_inst/buff[114][3] , \i11/fifo_inst/buff[114][4] , 
        \i11/fifo_inst/buff[114][5] , \i11/fifo_inst/buff[114][6] , \i11/fifo_inst/buff[114][7] , 
        \i11/fifo_inst/buff[115][0] , \i11/fifo_inst/buff[115][1] , \i11/fifo_inst/buff[115][2] , 
        \i11/fifo_inst/buff[115][3] , \i11/fifo_inst/buff[115][4] , \i11/fifo_inst/buff[115][5] , 
        \i11/fifo_inst/buff[115][6] , n1118, \i11/fifo_inst/buff[115][7] , 
        \i11/fifo_inst/buff[116][0] , \i11/fifo_inst/buff[116][1] , \i11/fifo_inst/buff[116][2] , 
        \i11/fifo_inst/buff[116][3] , n1124, \i11/fifo_inst/buff[116][4] , 
        n1126, n1127, \i11/fifo_inst/buff[116][5] , \i11/fifo_inst/buff[116][6] , 
        n1130, n1131, \i11/fifo_inst/buff[116][7] , n1133, \i11/fifo_inst/buff[117][0] , 
        \i11/fifo_inst/buff[117][1] , \i11/fifo_inst/buff[117][2] , \i11/fifo_inst/buff[117][3] , 
        \i11/fifo_inst/buff[117][4] , n1139, \i11/fifo_inst/buff[117][5] , 
        n1141, \i11/fifo_inst/buff[117][6] , \i11/fifo_inst/buff[117][7] , 
        \i11/fifo_inst/buff[118][0] , \i11/fifo_inst/buff[118][1] , \i11/fifo_inst/buff[118][2] , 
        \i11/fifo_inst/buff[118][3] , \i11/fifo_inst/buff[118][4] , \i11/fifo_inst/buff[118][5] , 
        n1150, \i11/fifo_inst/buff[118][6] , \i11/fifo_inst/buff[118][7] , 
        n1153, n1154, \i11/fifo_inst/buff[119][0] , n1156, n1157, 
        \i11/fifo_inst/buff[119][1] , n1159, n1160, \i11/fifo_inst/buff[119][2] , 
        \i11/fifo_inst/buff[119][3] , \i11/fifo_inst/buff[119][4] , \i11/fifo_inst/buff[119][5] , 
        \i11/fifo_inst/buff[119][6] , \i11/fifo_inst/buff[119][7] , n1167, 
        \i11/fifo_inst/buff[120][0] , n1169, n1170, \i11/fifo_inst/buff[120][1] , 
        n1172, n1173, \i11/fifo_inst/buff[120][2] , \i11/fifo_inst/buff[120][3] , 
        n1176, n1177, \i11/fifo_inst/buff[120][4] , n1179, n1180, 
        \i11/fifo_inst/buff[120][5] , n1182, n1183, \i11/fifo_inst/buff[120][6] , 
        \i11/fifo_inst/buff[120][7] , n1186, n1187, \i11/fifo_inst/buff[121][0] , 
        n1189, n1190, \i11/fifo_inst/buff[121][1] , n1192, n1193, 
        \i11/fifo_inst/buff[121][2] , \i11/fifo_inst/buff[121][3] , n1196, 
        n1197, \i11/fifo_inst/buff[121][4] , \i11/fifo_inst/buff[121][5] , 
        \i11/fifo_inst/buff[121][6] , \i11/fifo_inst/buff[121][7] , \i11/fifo_inst/buff[122][0] , 
        \i11/fifo_inst/buff[122][1] , \i11/fifo_inst/buff[122][2] , n1205, 
        n1206, \i11/fifo_inst/buff[122][3] , \i11/fifo_inst/buff[122][4] , 
        n1209, n1210, \i11/fifo_inst/buff[122][5] , \i11/fifo_inst/buff[122][6] , 
        \i11/fifo_inst/buff[122][7] , \i11/fifo_inst/buff[123][0] , \i11/fifo_inst/buff[123][1] , 
        \i11/fifo_inst/buff[123][2] , \i11/fifo_inst/buff[123][3] , \i11/fifo_inst/buff[123][4] , 
        n1219, n1220, \i11/fifo_inst/buff[123][5] , \i11/fifo_inst/buff[123][6] , 
        \i11/fifo_inst/buff[123][7] , n1224, n1225, \i11/fifo_inst/buff[124][0] , 
        \i11/fifo_inst/buff[124][1] , n1228, n1229, \i11/fifo_inst/buff[124][2] , 
        \i11/fifo_inst/buff[124][3] , n1232, n1233, \i11/fifo_inst/buff[124][4] , 
        \i11/fifo_inst/buff[124][5] , \i11/fifo_inst/buff[124][6] , n1237, 
        n1238, \i11/fifo_inst/buff[124][7] , \i11/fifo_inst/buff[125][0] , 
        n1241, n1242, \i11/fifo_inst/buff[125][1] , \i11/fifo_inst/buff[125][2] , 
        \i11/fifo_inst/buff[125][3] , \i11/fifo_inst/buff[125][4] , n1247, 
        n1248, \i11/fifo_inst/buff[125][5] , \i11/fifo_inst/buff[125][6] , 
        n1251, n1252, \i11/fifo_inst/buff[125][7] , n1254, n1255, 
        \i11/fifo_inst/buff[126][0] , \i11/fifo_inst/buff[126][1] , n1258, 
        n1259, \i11/fifo_inst/buff[126][2] , \i11/fifo_inst/buff[126][3] , 
        \i11/fifo_inst/buff[126][4] , \i11/fifo_inst/buff[126][5] , n1264, 
        \i11/fifo_inst/buff[126][6] , \i11/fifo_inst/buff[126][7] , n1267, 
        n1268, \i11/fifo_inst/buff[127][0] , \i11/fifo_inst/buff[127][1] , 
        \i11/fifo_inst/buff[127][2] , \i11/fifo_inst/buff[127][3] , n1273, 
        n1274, \i11/fifo_inst/buff[127][4] , \i11/fifo_inst/buff[127][5] , 
        n1277, n1278, \i11/fifo_inst/buff[127][6] , \i11/fifo_inst/buff[127][7] , 
        \spi_slave_inst/n95 , ceg_net5, \spi_slave_inst/n96 , \spi_slave_inst/n56 , 
        ceg_net37, \spi_slave_inst/n57 , \spi_slave_inst/sync_tx_en[0] , 
        \spi_slave_inst/n97 , tx_en, \spi_slave_inst/n58 , \spi_slave_inst/sync_mosi[0] , 
        \spi_slave_inst/n73 , ceg_net20, \spi_slave_inst/n98 , \spi_slave_inst/n139 , 
        ceg_net77, ceg_net98, \spi_slave_inst/n68 , ceg_net31, ceg_net34, 
        \spi_slave_inst/n54 , \spi_slave_inst/n55 , \spi_slave_inst/n138 , 
        \spi_slave_inst/n137 , \spi_slave_inst/n136 , \spi_slave_inst/n135 , 
        \spi_slave_inst/n134 , \spi_slave_inst/n133 , \spi_slave_inst/n132 , 
        \spi_slave_inst/n173 , \spi_slave_inst/n172 , \spi_slave_inst/n171 , 
        \spi_slave_inst/n170 , \spi_slave_inst/n169 , \spi_slave_inst/n168 , 
        \spi_slave_inst/n167 , \led_inst/n41 , \led_inst/n42 , \led_inst/n43 , 
        \led_inst/n44 , \led_inst/n45 , \led_inst/n48 , \led_inst/n46 , 
        \led_inst/n47 , \led_inst/n142 , \data_to_led[0] , rx_en_led, 
        \led_inst/LessThan_21/n48 , \led_inst/n141 , \led_inst/n140 , 
        \led_inst/n139 , \led_inst/n138 , \led_inst/n137 , \led_inst/n136 , 
        \led_inst/n135 , \led_inst/n134 , \led_inst/n133 , \led_inst/n132 , 
        \led_inst/n131 , \led_inst/n130 , \led_inst/n129 , \led_inst/n128 , 
        \led_inst/n127 , \led_inst/n126 , \led_inst/n125 , \led_inst/n124 , 
        \led_inst/n123 , \led_inst/n122 , \led_inst/n121 , \led_inst/n120 , 
        \led_inst/n119 , \data_to_led[1] , \data_to_led[2] , \data_to_led[3] , 
        \data_to_led[4] , \data_to_led[5] , \data_to_led[6] , \data_to_led[7] , 
        \data_to_fifo[5] , \i11/n128 , \data_to_gpo[0] , rx_en_gpo, 
        \data_to_fifo[4] , \data_to_gpo[1] , \data_to_gpo[2] , \data_to_gpo[3] , 
        \data_to_gpo[4] , \data_to_gpo[5] , \data_to_gpo[6] , \data_to_gpo[7] , 
        \data_to_fifo[0] , \i11/n130 , \data_to_fifo[3] , \data_to_fifo[7] , 
        \i11/n131 , \data_to_fifo[6] , \data_to_fifo[2] , \data_to_fifo[1] , 
        \i11/n129 , \tx_dac_fsm_inst/n68 , \tx_dac_fsm_inst/n42 , \tx_dac_fsm_inst/n344 , 
        n1410, n1411, \tx_dac_fsm_inst/n67 , \tx_dac_fsm_inst/n66 , 
        \tx_dac_fsm_inst/n65 , n1415, n1416, n1417, n1418, \tx_dac_fsm_inst/n258 , 
        \tx_dac_fsm_inst/n64 , \tx_dac_fsm_inst/n284 , data_to_dac, rx_en_dac, 
        \~tx_dac_fsm_inst/n431 , \~tx_dac_fsm_inst/n436 , \~tx_dac_fsm_inst/n441 , 
        n1436, n1437, n1438, n1439, \tx_dac_fsm_inst/n257 , \tx_dac_fsm_inst/n256 , 
        \tx_dac_fsm_inst/n255 , \tx_dac_fsm_inst/n254 , \tx_dac_fsm_inst/n253 , 
        \tx_dac_fsm_inst/n283 , \tx_dac_fsm_inst/n282 , \tx_dac_fsm_inst/n281 , 
        \tx_dac_fsm_inst/n280 , \tx_dac_fsm_inst/n279 , \fifo_inst/n153 , 
        ceg_net146, \fifo_inst/n162 , ceg_net164, \data_to_fifo_length[0] , 
        rx_en_fifo_length, rx_en_fifo, tx_en_fifo, \fifo_inst/n144 , 
        ceg_net242, \fifo_inst/n152 , \fifo_inst/n151 , \fifo_inst/n150 , 
        \fifo_inst/n149 , \fifo_inst/n148 , \fifo_inst/n147 , \fifo_inst/n146 , 
        \fifo_inst/n161 , \fifo_inst/n160 , \fifo_inst/n159 , \fifo_inst/n158 , 
        \fifo_inst/n157 , \fifo_inst/n156 , \fifo_inst/n155 , \data_to_fifo_length[1] , 
        \data_to_fifo_length[2] , \data_to_fifo_length[3] , \data_to_fifo_length[4] , 
        \data_to_fifo_length[5] , \data_to_fifo_length[6] , \data_to_fifo_length[7] , 
        \i11/n132 , \fifo_inst/n143 , \fifo_inst/n142 , \fifo_inst/n141 , 
        \fifo_inst/n140 , \fifo_inst/n139 , \fifo_inst/n138 , \fifo_inst/n137 , 
        \i11/n127 , \i11/n126 , \i11/n125 , \i11/n124 , \i11/n123 , 
        \i11/n122 , \i11/n121 , \i11/n120 , \i11/n119 , \i11/n118 , 
        \i11/n117 , \i11/n116 , \i11/n115 , \i11/n114 , \i11/n113 , 
        \i11/n112 , \i11/n111 , \i11/n110 , \i11/n109 , \i11/n108 , 
        \i11/n107 , \i11/n106 , \i11/n105 , \i11/n104 , \i11/n103 , 
        \i11/n102 , \i11/n101 , \i11/n100 , \i11/n99 , \i11/n98 , 
        \i11/n97 , \i11/n96 , \i11/n95 , \i11/n94 , \i11/n93 , \i11/n92 , 
        \i11/n91 , \i11/n90 , \i11/n89 , \i11/n88 , \i11/n87 , \i11/n86 , 
        \i11/n85 , \i11/n84 , \i11/n83 , \i11/n82 , \i11/n81 , \i11/n80 , 
        \i11/n79 , \i11/n78 , \i11/n77 , \i11/n76 , \i11/n75 , \i11/n74 , 
        \i11/n73 , \i11/n72 , \i11/n71 , \i11/n70 , \i11/n69 , \i11/n68 , 
        \i11/n67 , \i11/n66 , \i11/n65 , \i11/n64 , \i11/n63 , \i11/n62 , 
        \i11/n61 , \i11/n60 , \i11/n59 , \i11/n58 , \i11/n57 , \i11/n56 , 
        \i11/n55 , \i11/n54 , \i11/n53 , \i11/n52 , \i11/n51 , \i11/n50 , 
        \i11/n49 , \i11/n48 , \i11/n47 , \i11/n46 , \i11/n45 , \i11/n44 , 
        \i11/n43 , \i11/n42 , \i11/n41 , \i11/n40 , \i11/n39 , \i11/n38 , 
        \i11/n37 , \i11/n36 , \i11/n35 , \i11/n34 , \i11/n33 , \i11/n32 , 
        \i11/n31 , \i11/n30 , \i11/n29 , \i11/n28 , \i11/n27 , \i11/n26 , 
        \i11/n25 , \i11/n24 , \i11/n23 , \i11/n22 , \i11/n21 , \i11/n20 , 
        \i11/n19 , n1617, \i11/n18 , \i11/n17 , \i11/n16 , n1628, 
        \i11/n15 , n1633, \i11/n14 , \i11/n13 , \i11/n12 , \i11/n11 , 
        \i11/n10 , \i11/n9 , \i11/n8 , \i11/n7 , \i11/n6 , \tx_slowclk~O , 
        \pll_clk~O , n2612, n2611, n2610, n2609, \i11/n5 , n2608, 
        \tx_dac_fsm_inst/dctr[4]~FF_frt_0_q_pinv , \tx_dac_fsm_inst/dctr[1]~FF_frt_1_q , 
        \tx_dac_fsm_inst/dctr[4]~FF_frt_0_q , n1703, n1704, n1705, n1706, 
        n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, 
        n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
        n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, 
        n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, 
        n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
        n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, 
        n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
        n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, 
        n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, 
        n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
        n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, 
        n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, 
        n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, 
        n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, 
        n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
        n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, 
        n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
        n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, 
        n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, 
        n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
        n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, 
        n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
        n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, 
        n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, 
        n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
        n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, 
        n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
        n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, 
        n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, 
        n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
        n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, 
        n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
        n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, 
        n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, 
        n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
        n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, 
        n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
        n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, 
        n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, 
        n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
        n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, 
        n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
        n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, 
        n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, 
        n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
        n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, 
        n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
        n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, 
        n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, 
        n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
        n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, 
        n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
        n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, 
        n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, 
        n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
        n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, 
        n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
        n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, 
        n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, 
        n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, 
        n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, 
        n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
        n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, 
        n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, 
        n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
        n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, 
        n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
        n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, 
        n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, 
        n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, 
        n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, 
        n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
        n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, 
        n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, 
        n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, 
        n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, 
        n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
        n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, 
        n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, 
        n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, 
        n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, 
        n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
        n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, 
        n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, 
        n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, 
        n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, 
        n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
        n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, 
        n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, 
        n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
        n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, 
        n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, 
        n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, 
        n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, 
        n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, 
        n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, 
        n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, 
        n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
        n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, 
        n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, 
        n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, 
        n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, 
        n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, 
        n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, 
        n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
        n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, 
        n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, 
        n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, 
        n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, 
        n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, 
        n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, 
        n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, 
        n2603, n2604, n2605, n2606, n2607;
    
    EFX_LUT4 \tx_dac_fsm_inst/dlatchrs_162/i1  (.I0(n1410), .I1(n125), .I2(n1411), 
            .O(n125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/dlatchrs_162/i1 .LUTMASK = 16'hacac;
    EFX_LUT4 \tx_dac_fsm_inst/i116  (.I0(n1415), .I1(n130), .I2(n1416), 
            .O(n130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/i116 .LUTMASK = 16'hacac;
    EFX_FF \reg_addr[3]~FF  (.D(\spi_slave_inst/n95 ), .CE(ceg_net5), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\reg_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(114)
    defparam \reg_addr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \reg_addr[3]~FF .CE_POLARITY = 1'b0;
    defparam \reg_addr[3]~FF .SR_POLARITY = 1'b0;
    defparam \reg_addr[3]~FF .D_POLARITY = 1'b1;
    defparam \reg_addr[3]~FF .SR_SYNC = 1'b0;
    defparam \reg_addr[3]~FF .SR_VALUE = 1'b0;
    defparam \reg_addr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \reg_addr[2]~FF  (.D(\spi_slave_inst/n96 ), .CE(ceg_net5), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\reg_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(114)
    defparam \reg_addr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \reg_addr[2]~FF .CE_POLARITY = 1'b0;
    defparam \reg_addr[2]~FF .SR_POLARITY = 1'b0;
    defparam \reg_addr[2]~FF .D_POLARITY = 1'b1;
    defparam \reg_addr[2]~FF .SR_SYNC = 1'b0;
    defparam \reg_addr[2]~FF .SR_VALUE = 1'b0;
    defparam \reg_addr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/bitcnt[2]~FF  (.D(\spi_slave_inst/n56 ), .CE(ceg_net37), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/bitcnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/bitcnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[2]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[2]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/bitcnt[2]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/bitcnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/bitcnt[1]~FF  (.D(\spi_slave_inst/n57 ), .CE(ceg_net37), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/bitcnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/bitcnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[1]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[1]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/bitcnt[1]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/bitcnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_tx_en[1]~FF  (.D(\spi_slave_inst/sync_tx_en[0] ), 
           .CE(1'b1), .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/sync_tx_en[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_tx_en[1]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_tx_en[1]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_tx_en[1]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_tx_en[1]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_tx_en[1]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_tx_en[1]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/sync_tx_en[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \reg_addr[1]~FF  (.D(\spi_slave_inst/n97 ), .CE(ceg_net5), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\reg_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(114)
    defparam \reg_addr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \reg_addr[1]~FF .CE_POLARITY = 1'b0;
    defparam \reg_addr[1]~FF .SR_POLARITY = 1'b0;
    defparam \reg_addr[1]~FF .D_POLARITY = 1'b1;
    defparam \reg_addr[1]~FF .SR_SYNC = 1'b0;
    defparam \reg_addr[1]~FF .SR_VALUE = 1'b0;
    defparam \reg_addr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_tx_en[0]_2~FF  (.D(tx_en), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\spi_slave_inst/sync_tx_en[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_tx_en[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_tx_en[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_tx_en[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_tx_en[0]_2~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_tx_en[0]_2~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_tx_en[0]_2~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/sync_tx_en[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/bitcnt[0]~FF  (.D(\spi_slave_inst/n58 ), .CE(ceg_net37), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/bitcnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/bitcnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[0]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[0]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/bitcnt[0]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/bitcnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_mosi[1]~FF  (.D(\spi_slave_inst/sync_mosi[0] ), 
           .CE(1'b1), .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/sync_mosi[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_mosi[1]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_mosi[1]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_mosi[1]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_mosi[1]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_mosi[1]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_mosi[1]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/sync_mosi[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rw_out~FF  (.D(\spi_slave_inst/n73 ), .CE(ceg_net20), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(rw_out)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(103)
    defparam \rw_out~FF .CLK_POLARITY = 1'b1;
    defparam \rw_out~FF .CE_POLARITY = 1'b0;
    defparam \rw_out~FF .SR_POLARITY = 1'b0;
    defparam \rw_out~FF .D_POLARITY = 1'b1;
    defparam \rw_out~FF .SR_SYNC = 1'b0;
    defparam \rw_out~FF .SR_VALUE = 1'b0;
    defparam \rw_out~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \reg_addr[0]~FF  (.D(\spi_slave_inst/n98 ), .CE(ceg_net5), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\reg_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(114)
    defparam \reg_addr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \reg_addr[0]~FF .CE_POLARITY = 1'b0;
    defparam \reg_addr[0]~FF .SR_POLARITY = 1'b0;
    defparam \reg_addr[0]~FF .D_POLARITY = 1'b1;
    defparam \reg_addr[0]~FF .SR_SYNC = 1'b0;
    defparam \reg_addr[0]~FF .SR_VALUE = 1'b0;
    defparam \reg_addr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[0]~FF  (.D(\spi_slave_inst/n139 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[0]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[0]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[0]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[0]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[0]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[0]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[0]~FF  (.D(\spi_slave_inst/n98 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[0]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[0]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[0]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[0]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[0]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[0]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \addr_dv~FF  (.D(\spi_slave_inst/n68 ), .CE(ceg_net31), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(addr_dv)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(155)
    defparam \addr_dv~FF .CLK_POLARITY = 1'b1;
    defparam \addr_dv~FF .CE_POLARITY = 1'b0;
    defparam \addr_dv~FF .SR_POLARITY = 1'b0;
    defparam \addr_dv~FF .D_POLARITY = 1'b0;
    defparam \addr_dv~FF .SR_SYNC = 1'b0;
    defparam \addr_dv~FF .SR_VALUE = 1'b0;
    defparam \addr_dv~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rxdv~FF  (.D(\spi_slave_inst/n68 ), .CE(ceg_net34), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(rxdv)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(165)
    defparam \rxdv~FF .CLK_POLARITY = 1'b1;
    defparam \rxdv~FF .CE_POLARITY = 1'b0;
    defparam \rxdv~FF .SR_POLARITY = 1'b0;
    defparam \rxdv~FF .D_POLARITY = 1'b0;
    defparam \rxdv~FF .SR_SYNC = 1'b0;
    defparam \rxdv~FF .SR_VALUE = 1'b0;
    defparam \rxdv~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_sclk[0]~FF  (.D(SCLK), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\spi_slave_inst/sync_sclk[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_sclk[0]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[0]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[0]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_sclk[0]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[0]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_sclk[0]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/sync_sclk[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/bitcnt[4]~FF  (.D(\spi_slave_inst/n54 ), .CE(ceg_net37), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/bitcnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/bitcnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[4]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[4]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/bitcnt[4]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/bitcnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/bitcnt[3]~FF  (.D(\spi_slave_inst/n55 ), .CE(ceg_net37), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/bitcnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/bitcnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[3]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[3]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/bitcnt[3]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/bitcnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_mosi[0]_2~FF  (.D(MOSI), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\spi_slave_inst/sync_mosi[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_mosi[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_mosi[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_mosi[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_mosi[0]_2~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_mosi[0]_2~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_mosi[0]_2~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/sync_mosi[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_ss[0]~FF  (.D(SSB), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\spi_slave_inst/sync_ss[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_ss[0]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[0]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[0]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_ss[0]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[0]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_ss[0]~FF .SR_VALUE = 1'b1;
    defparam \spi_slave_inst/sync_ss[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[1]~FF  (.D(\spi_slave_inst/n138 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[1]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[1]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[1]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[1]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[1]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[2]~FF  (.D(\spi_slave_inst/n137 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[2]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[2]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[2]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[2]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[2]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[2]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[3]~FF  (.D(\spi_slave_inst/n136 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[3]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[3]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[3]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[3]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[3]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[3]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[4]~FF  (.D(\spi_slave_inst/n135 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[4]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[4]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[4]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[4]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[4]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[4]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[5]~FF  (.D(\spi_slave_inst/n134 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[5]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[5]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[5]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[5]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[5]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[5]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[6]~FF  (.D(\spi_slave_inst/n133 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[6]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[6]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[6]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[6]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[6]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[6]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[7]~FF  (.D(\spi_slave_inst/n132 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[7]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[7]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[7]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[7]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[7]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[7]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[1]~FF  (.D(\spi_slave_inst/n173 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[1]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[1]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[1]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[1]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[1]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[1]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[2]~FF  (.D(\spi_slave_inst/n172 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[2]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[2]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[2]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[2]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[2]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[2]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[3]~FF  (.D(\spi_slave_inst/n171 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[3]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[3]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[3]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[3]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[3]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[3]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[4]~FF  (.D(\spi_slave_inst/n170 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[4]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[4]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[4]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[4]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[4]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[4]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[5]~FF  (.D(\spi_slave_inst/n169 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[5]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[5]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[5]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[5]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[5]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[5]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[6]~FF  (.D(\spi_slave_inst/n168 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[6]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[6]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[6]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[6]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[6]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[6]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[7]~FF  (.D(\spi_slave_inst/n167 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[7]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[7]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[7]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[7]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[7]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[7]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_sclk[1]~FF  (.D(\spi_slave_inst/sync_sclk[0] ), 
           .CE(1'b1), .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/sync_sclk[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_sclk[1]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[1]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[1]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_sclk[1]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[1]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_sclk[1]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/sync_sclk[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_sclk[2]~FF  (.D(\spi_slave_inst/sync_sclk[1] ), 
           .CE(1'b1), .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/sync_sclk[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_sclk[2]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[2]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[2]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_sclk[2]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[2]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_sclk[2]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/sync_sclk[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_ss[1]~FF  (.D(\spi_slave_inst/sync_ss[0] ), 
           .CE(1'b1), .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/sync_ss[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_ss[1]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[1]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[1]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_ss[1]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[1]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_ss[1]~FF .SR_VALUE = 1'b1;
    defparam \spi_slave_inst/sync_ss[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_ss[2]~FF  (.D(\spi_slave_inst/sync_ss[1] ), 
           .CE(1'b1), .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/sync_ss[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_ss[2]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[2]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[2]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_ss[2]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[2]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_ss[2]~FF .SR_VALUE = 1'b1;
    defparam \spi_slave_inst/sync_ss[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[7]~FF  (.D(\led_inst/n41 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[7]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[7]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[7]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[7]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[7]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[7]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[6]~FF  (.D(\led_inst/n42 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[6]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[6]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[6]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[6]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[6]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[6]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[5]~FF  (.D(\led_inst/n43 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[5]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[5]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[5]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[5]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[5]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[5]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[4]~FF  (.D(\led_inst/n44 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[4]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[4]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[4]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[4]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[4]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[4]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[3]~FF  (.D(\led_inst/n45 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[3]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[3]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[3]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[3]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[3]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[3]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[0]~FF  (.D(\led_inst/n48 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[0]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[0]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[0]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[0]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[0]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[0]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[2]~FF  (.D(\led_inst/n46 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[2]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[2]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[2]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[2]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[2]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[2]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[1]~FF  (.D(\led_inst/n47 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[1]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[1]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[1]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[1]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[1]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[1]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[0]~FF  (.D(\led_inst/n142 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[0]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[0]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[0]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[0]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[0]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[0]~FF  (.D(\data_to_led[0] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[0]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[0]~FF .SR_VALUE = 1'b1;
    defparam \led_inst/ctr_cfg_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led0~FF  (.D(led0), .CE(\led_inst/LessThan_21/n48 ), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(led0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led0~FF .CLK_POLARITY = 1'b1;
    defparam \led0~FF .CE_POLARITY = 1'b1;
    defparam \led0~FF .SR_POLARITY = 1'b0;
    defparam \led0~FF .D_POLARITY = 1'b0;
    defparam \led0~FF .SR_SYNC = 1'b0;
    defparam \led0~FF .SR_VALUE = 1'b0;
    defparam \led0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led1~FF  (.D(led0), .CE(\led_inst/LessThan_21/n48 ), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(led1)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led1~FF .CLK_POLARITY = 1'b1;
    defparam \led1~FF .CE_POLARITY = 1'b1;
    defparam \led1~FF .SR_POLARITY = 1'b0;
    defparam \led1~FF .D_POLARITY = 1'b1;
    defparam \led1~FF .SR_SYNC = 1'b0;
    defparam \led1~FF .SR_VALUE = 1'b1;
    defparam \led1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[1]~FF  (.D(\led_inst/n141 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[1]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[1]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[1]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[1]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[2]~FF  (.D(\led_inst/n140 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[2]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[2]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[2]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[2]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[3]~FF  (.D(\led_inst/n139 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[3]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[3]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[3]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[3]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[4]~FF  (.D(\led_inst/n138 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[4]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[4]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[4]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[4]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[5]~FF  (.D(\led_inst/n137 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[5]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[5]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[5]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[5]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[6]~FF  (.D(\led_inst/n136 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[6]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[6]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[6]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[6]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[6]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[7]~FF  (.D(\led_inst/n135 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[7]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[7]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[7]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[7]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[7]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[8]~FF  (.D(\led_inst/n134 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[8]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[8]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[8]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[8]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[8]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[9]~FF  (.D(\led_inst/n133 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[9]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[9]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[9]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[9]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[9]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[10]~FF  (.D(\led_inst/n132 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[10]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[10]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[10]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[10]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[10]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[11]~FF  (.D(\led_inst/n131 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[11]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[11]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[11]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[11]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[11]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[12]~FF  (.D(\led_inst/n130 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[12]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[12]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[12]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[12]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[12]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[13]~FF  (.D(\led_inst/n129 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[13]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[13]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[13]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[13]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[13]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[14]~FF  (.D(\led_inst/n128 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[14]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[14]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[14]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[14]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[14]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[15]~FF  (.D(\led_inst/n127 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[15]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[15]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[15]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[15]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[15]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[16]~FF  (.D(\led_inst/n126 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[16]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[16]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[16]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[16]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[16]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[16]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[17]~FF  (.D(\led_inst/n125 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[17]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[17]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[17]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[17]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[17]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[17]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[18]~FF  (.D(\led_inst/n124 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[18]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[18]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[18]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[18]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[18]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[18]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[19]~FF  (.D(\led_inst/n123 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[19]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[19]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[19]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[19]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[19]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[19]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[20]~FF  (.D(\led_inst/n122 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[20]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[20]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[20]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[20]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[20]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[20]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[21]~FF  (.D(\led_inst/n121 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[21]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[21]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[21]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[21]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[21]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[21]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[22]~FF  (.D(\led_inst/n120 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[22]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[22]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[22]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[22]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[22]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[22]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[23]~FF  (.D(\led_inst/n119 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[23]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[23]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[23]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[23]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[23]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[23]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[1]~FF  (.D(\data_to_led[1] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[1]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/ctr_cfg_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[2]~FF  (.D(\data_to_led[2] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[2]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[2]~FF .SR_VALUE = 1'b1;
    defparam \led_inst/ctr_cfg_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[3]~FF  (.D(\data_to_led[3] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[3]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[3]~FF .SR_VALUE = 1'b1;
    defparam \led_inst/ctr_cfg_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[4]~FF  (.D(\data_to_led[4] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[4]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[4]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[4]~FF .SR_VALUE = 1'b1;
    defparam \led_inst/ctr_cfg_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[5]~FF  (.D(\data_to_led[5] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[5]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[5]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/ctr_cfg_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[6]~FF  (.D(\data_to_led[6] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[6]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[6]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[6]~FF .SR_VALUE = 1'b1;
    defparam \led_inst/ctr_cfg_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[7]~FF  (.D(\data_to_led[7] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[7]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[7]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/ctr_cfg_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[4][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[4][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[4][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[4][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[4][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[0]~FF  (.D(\data_to_gpo[0] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[0]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[4][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[4][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[4][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[4][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[4][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[1]~FF  (.D(\data_to_gpo[1] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[1]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[2]~FF  (.D(\data_to_gpo[2] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[2]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[3]~FF  (.D(\data_to_gpo[3] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[3]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[4]~FF  (.D(\data_to_gpo[4] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[4]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[4]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[5]~FF  (.D(\data_to_gpo[5] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[5]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[5]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[6]~FF  (.D(\data_to_gpo[6] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[6]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[6]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[7]~FF  (.D(\data_to_gpo[7] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[7]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[7]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[2][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[2][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[2][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[2][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[2][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[2][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[2][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[2][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[2][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[2][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[1][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[1][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[1][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[1][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[1][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[1][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[1][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[1][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[1][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[1][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[1][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[1][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[1][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[1][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[1][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[2][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[2][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[2][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[2][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[2][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[4][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[4][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[4][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[4][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[4][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[2][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[2][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[2][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[2][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[2][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[4][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[4][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[4][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[4][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[4][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[1][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[1][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[1][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[1][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[1][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[4][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[4][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[4][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[4][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[4][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[4][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[4][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[4][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[4][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[4][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[3][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[3][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[3][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[3][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[3][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[3][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[3][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[3][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[3][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[3][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[3][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[3][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[3][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[3][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[3][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[3][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[3][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[3][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[3][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[3][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[3][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[3][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[3][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[3][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[3][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[3][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[3][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[3][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[3][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[3][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[3][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[3][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[3][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[3][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[3][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[3][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[3][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[3][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[3][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[3][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[3][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[2][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[2][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[2][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[2][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[2][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_ctr[0]~FF  (.D(\tx_dac_fsm_inst/n68 ), .CE(\tx_dac_fsm_inst/n42 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_ctr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_ctr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_pos[0]~FF  (.D(\tx_dac_fsm_inst/sym_pos[0] ), 
           .CE(\tx_dac_fsm_inst/n344 ), .CLK(\tx_slowclk~O ), .SR(reset_n), 
           .Q(\tx_dac_fsm_inst/sym_pos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_pos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[0]~FF .D_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/state_reg[0]~FF  (.D(n125), .CE(1'b1), .CLK(\tx_slowclk~O ), 
           .SR(reset_n), .Q(\tx_dac_fsm_inst/state_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(113)
    defparam \tx_dac_fsm_inst/state_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_ctr[1]~FF  (.D(\tx_dac_fsm_inst/n67 ), .CE(\tx_dac_fsm_inst/n42 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_ctr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_ctr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[1]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_ctr[2]~FF  (.D(\tx_dac_fsm_inst/n66 ), .CE(\tx_dac_fsm_inst/n42 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_ctr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_ctr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[2]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[2]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[2]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[2]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[2]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_ctr[3]~FF  (.D(\tx_dac_fsm_inst/n65 ), .CE(\tx_dac_fsm_inst/n42 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_ctr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_ctr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[3]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[3]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[3]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[3]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[3]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[2][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[2][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[2][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[2][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[2][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[2][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[2][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[2][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[2][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[2][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/zctr[0]~FF  (.D(\tx_dac_fsm_inst/n258 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/zctr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(200)
    defparam \tx_dac_fsm_inst/zctr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_ctr[4]~FF  (.D(\tx_dac_fsm_inst/n64 ), .CE(\tx_dac_fsm_inst/n42 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_ctr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_ctr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[4]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[4]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[4]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[4]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[4]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dctr[0]~FF  (.D(\tx_dac_fsm_inst/n284 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/dctr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(211)
    defparam \tx_dac_fsm_inst/dctr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dac_config_reg[0]~FF  (.D(data_to_dac), .CE(rx_en_dac), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/dac_config_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(51)
    defparam \tx_dac_fsm_inst/dac_config_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dac_config_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dac_config_reg[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dac_config_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dac_config_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dac_config_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dac_config_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_pos[1]~FF  (.D(\~tx_dac_fsm_inst/n431 ), .CE(\tx_dac_fsm_inst/n344 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_pos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_pos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[1]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_pos[2]~FF  (.D(\~tx_dac_fsm_inst/n436 ), .CE(\tx_dac_fsm_inst/n344 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_pos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_pos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[2]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[2]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[2]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[2]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[2]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_pos[3]~FF  (.D(\~tx_dac_fsm_inst/n441 ), .CE(\tx_dac_fsm_inst/n344 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_pos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_pos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[3]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[3]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[3]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[3]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[3]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/state_reg[1]~FF  (.D(n150), .CE(1'b1), .CLK(\tx_slowclk~O ), 
           .SR(reset_n), .Q(\tx_dac_fsm_inst/state_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(113)
    defparam \tx_dac_fsm_inst/state_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/state_reg[2]~FF  (.D(n151), .CE(1'b1), .CLK(\tx_slowclk~O ), 
           .SR(reset_n), .Q(\tx_dac_fsm_inst/state_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(113)
    defparam \tx_dac_fsm_inst/state_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[2]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/state_reg[3]~FF  (.D(n152), .CE(1'b1), .CLK(\tx_slowclk~O ), 
           .SR(reset_n), .Q(\tx_dac_fsm_inst/state_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(113)
    defparam \tx_dac_fsm_inst/state_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[3]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/zctr[1]~FF  (.D(\tx_dac_fsm_inst/n257 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/zctr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(200)
    defparam \tx_dac_fsm_inst/zctr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[1]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/zctr[2]~FF  (.D(\tx_dac_fsm_inst/n256 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/zctr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(200)
    defparam \tx_dac_fsm_inst/zctr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[2]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[2]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[2]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[2]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[2]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/zctr[3]~FF  (.D(\tx_dac_fsm_inst/n255 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/zctr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(200)
    defparam \tx_dac_fsm_inst/zctr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[3]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[3]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[3]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[3]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[3]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/zctr[4]~FF  (.D(\tx_dac_fsm_inst/n254 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/zctr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(200)
    defparam \tx_dac_fsm_inst/zctr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[4]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[4]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[4]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[4]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[4]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/zctr[5]~FF  (.D(\tx_dac_fsm_inst/n253 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/zctr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(200)
    defparam \tx_dac_fsm_inst/zctr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[5]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[5]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[5]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[5]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[5]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dctr[1]~FF  (.D(\tx_dac_fsm_inst/n283 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/dctr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(211)
    defparam \tx_dac_fsm_inst/dctr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[1]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dctr[2]~FF  (.D(\tx_dac_fsm_inst/n282 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/dctr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(211)
    defparam \tx_dac_fsm_inst/dctr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[2]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[2]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[2]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[2]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[2]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dctr[3]~FF  (.D(\tx_dac_fsm_inst/n281 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/dctr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(211)
    defparam \tx_dac_fsm_inst/dctr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[3]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[3]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[3]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[3]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[3]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dctr[4]~FF  (.D(\tx_dac_fsm_inst/n280 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/dctr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(211)
    defparam \tx_dac_fsm_inst/dctr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[4]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[4]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[4]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[4]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[4]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dctr[5]~FF  (.D(\tx_dac_fsm_inst/n279 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/dctr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(211)
    defparam \tx_dac_fsm_inst/dctr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[5]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[5]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[5]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[5]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[5]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[0]~FF  (.D(\fifo_inst/n153 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/wr_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[0]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[0]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[0]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[0]~FF  (.D(\fifo_inst/n162 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/rd_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[0]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[0]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[0]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[0]~FF  (.D(\data_to_fifo_length[0] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/length[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[0]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[0]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[0]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[0]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[0]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/sync_wr[0]~FF  (.D(rx_en_fifo), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\fifo_inst/sync_wr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/sync_wr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/sync_wr[0]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/sync_wr[0]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/sync_wr[0]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/sync_wr[0]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/sync_wr[0]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/sync_wr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/sync_rd[0]~FF  (.D(tx_en_fifo), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\fifo_inst/sync_rd[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/sync_rd[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/sync_rd[0]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/sync_rd[0]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/sync_rd[0]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/sync_rd[0]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/sync_rd[0]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/sync_rd[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[0]~FF  (.D(\fifo_inst/n144 ), .CE(ceg_net242), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/buff_head[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[0]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[0]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[0]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[0]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[0]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[1]~FF  (.D(\fifo_inst/n152 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/wr_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[1]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[1]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[1]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[2]~FF  (.D(\fifo_inst/n151 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/wr_index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[2]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[2]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[2]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[2]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[2]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[3]~FF  (.D(\fifo_inst/n150 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/wr_index[3]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[3]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[3]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[3]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[3]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[3]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[4]~FF  (.D(\fifo_inst/n149 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/wr_index[4]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[4]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[4]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[4]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[4]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[4]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[5]~FF  (.D(\fifo_inst/n148 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/wr_index[5]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[5]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[5]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[5]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[5]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[5]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[6]~FF  (.D(\fifo_inst/n147 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/wr_index[6]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[6]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[6]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[6]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[6]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[6]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[7]~FF  (.D(\fifo_inst/n146 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/wr_index[7]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[7]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[7]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[7]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[7]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[7]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[1]~FF  (.D(\fifo_inst/n161 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/rd_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[1]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[1]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[1]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[2]~FF  (.D(\fifo_inst/n160 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/rd_index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[2]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[2]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[2]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[2]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[2]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[3]~FF  (.D(\fifo_inst/n159 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/rd_index[3]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[3]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[3]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[3]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[3]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[3]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[4]~FF  (.D(\fifo_inst/n158 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/rd_index[4]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[4]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[4]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[4]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[4]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[4]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[5]~FF  (.D(\fifo_inst/n157 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/rd_index[5]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[5]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[5]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[5]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[5]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[5]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[6]~FF  (.D(\fifo_inst/n156 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/rd_index[6]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[6]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[6]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[6]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[6]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[6]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[7]~FF  (.D(\fifo_inst/n155 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/rd_index[7]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[7]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[7]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[7]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[7]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[7]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[1]~FF  (.D(\data_to_fifo_length[1] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/length[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[1]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[1]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[1]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[1]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[1]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[2]~FF  (.D(\data_to_fifo_length[2] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/length[2]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[2]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[2]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[2]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[2]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[2]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[3]~FF  (.D(\data_to_fifo_length[3] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/length[3]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[3]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[3]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[3]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[3]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[3]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[4]~FF  (.D(\data_to_fifo_length[4] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/length[4]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[4]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[4]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[4]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[4]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[4]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[5]~FF  (.D(\data_to_fifo_length[5] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/length[5]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[5]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[5]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[5]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[5]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[5]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[6]~FF  (.D(\data_to_fifo_length[6] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/length[6]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[6]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[6]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[6]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[6]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[6]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[7]~FF  (.D(\data_to_fifo_length[7] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/length[7]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[7]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[7]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[7]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[7]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[7]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/sync_wr[1]~FF  (.D(\fifo_inst/sync_wr[0] ), .CE(1'b1), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/sync_wr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/sync_wr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/sync_wr[1]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/sync_wr[1]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/sync_wr[1]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/sync_wr[1]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/sync_wr[1]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/sync_wr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/sync_rd[1]~FF  (.D(\fifo_inst/sync_rd[0] ), .CE(1'b1), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/sync_rd[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/sync_rd[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/sync_rd[1]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/sync_rd[1]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/sync_rd[1]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/sync_rd[1]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/sync_rd[1]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/sync_rd[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[0][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[0][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[0][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[0][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[0][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[0][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[0][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[0][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[1][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[1][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[1][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[1][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[1][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[1][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[1][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[1][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[1][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[1][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[2][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[2][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[2][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[2][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[2][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[2][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[0][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[0][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[0][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[0][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[0][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[0][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[0][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[0][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[0][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[1][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[1][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[1][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[1][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[1][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[1][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[1][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[1][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[1][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[1][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[1][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[1]~FF  (.D(\fifo_inst/n143 ), .CE(ceg_net242), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/buff_head[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[1]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[1]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[1]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[1]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[1]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[2]~FF  (.D(\fifo_inst/n142 ), .CE(ceg_net242), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/buff_head[2]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[2]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[2]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[2]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[2]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[2]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[3]~FF  (.D(\fifo_inst/n141 ), .CE(ceg_net242), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/buff_head[3]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[3]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[3]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[3]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[3]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[3]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[4]~FF  (.D(\fifo_inst/n140 ), .CE(ceg_net242), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/buff_head[4]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[4]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[4]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[4]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[4]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[4]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[5]~FF  (.D(\fifo_inst/n139 ), .CE(ceg_net242), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/buff_head[5]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[5]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[5]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[5]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[5]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[5]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[6]~FF  (.D(\fifo_inst/n138 ), .CE(ceg_net242), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/buff_head[6]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[6]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[6]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[6]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[6]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[6]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[7]~FF  (.D(\fifo_inst/n137 ), .CE(ceg_net242), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(84)
    defparam \fifo_inst/buff_head[7]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[7]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[7]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[7]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[7]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[7]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[4][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[4][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[4][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[4][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[4][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[4][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[4][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[4][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[4][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[4][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[4][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[5][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[5][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[5][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[5][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[5][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[5][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[5][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[5][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[5][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[5][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[5][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[5][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[5][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[5][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[5][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[5][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[5][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[5][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[5][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[5][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[5][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[5][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[5][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[5][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[5][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[5][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[5][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[5][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[5][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[5][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[5][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[5][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[5][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[5][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[5][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[5][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[5][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[5][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[5][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[5][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[5][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[6][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[6][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[6][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[6][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[6][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[6][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[6][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[6][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[6][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[6][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[6][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[6][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[6][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[6][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[6][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[6][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[6][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[6][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[6][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[6][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[6][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[6][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[6][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[6][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[6][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[6][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[6][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[6][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[6][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[6][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[6][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[6][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[6][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[6][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[6][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[6][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[6][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[6][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[6][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[6][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[6][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[7][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[7][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[7][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[7][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[7][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[7][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[7][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[7][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[7][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[7][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[7][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[7][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[7][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[7][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[7][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[7][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[7][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[7][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[7][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[7][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[7][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[7][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[7][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[7][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[7][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[7][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[7][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[7][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[7][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[7][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[7][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[7][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[7][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[7][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[7][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[7][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[7][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[7][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[7][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[7][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[7][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[8][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[8][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[8][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[8][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[8][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[8][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[8][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[8][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[8][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[8][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[8][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[8][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[8][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[8][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[8][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[8][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[8][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[8][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[8][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[8][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[8][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[8][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[8][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[8][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[8][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[8][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[8][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[8][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[8][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[8][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[8][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[8][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[8][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[8][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[8][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[8][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[8][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[8][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[8][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[8][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[8][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[9][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[9][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[9][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[9][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[9][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[9][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[9][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[9][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[9][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[9][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[9][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[9][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[9][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[9][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[9][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[9][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[9][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[9][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[9][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[9][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[9][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[9][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[9][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[9][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[9][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[9][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[9][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[9][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[9][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[9][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[9][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[9][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[9][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[9][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[9][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[9][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[9][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[9][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[9][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[9][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[9][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[10][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[10][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[10][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[10][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[10][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[10][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[10][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[10][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[10][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[10][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[10][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[10][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[10][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[10][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[10][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[10][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[10][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[10][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[10][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[10][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[10][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[10][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[10][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[10][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[10][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[10][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[10][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[10][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[10][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[10][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[10][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[10][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[10][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[10][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[10][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[10][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[10][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[10][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[10][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[10][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[10][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[11][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[11][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[11][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[11][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[11][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[11][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[11][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[11][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[11][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[11][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[11][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[11][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[11][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[11][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[11][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[11][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[11][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[11][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[11][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[11][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[11][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[11][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[11][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[11][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[11][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[11][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[11][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[11][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[11][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[11][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[11][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[11][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[11][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[11][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[11][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[11][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[11][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[11][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[11][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[11][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[11][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[12][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[12][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[12][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[12][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[12][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[12][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[12][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[12][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[12][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[12][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[12][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[12][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[12][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[12][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[12][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[12][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[12][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[12][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[12][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[12][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[12][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[12][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[12][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[12][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[12][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[12][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[12][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[12][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[12][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[12][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[12][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[12][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[12][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[12][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[12][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[12][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[12][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[12][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[12][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[12][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[12][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[13][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[13][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[13][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[13][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[13][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[13][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[13][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[13][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[13][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[13][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[13][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[13][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[13][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[13][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[13][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[13][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[13][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[13][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[13][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[13][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[13][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[13][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[13][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[13][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[13][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[13][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[13][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[13][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[13][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[13][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[13][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[13][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[13][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[13][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[13][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[13][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[13][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[13][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[13][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[13][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[13][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[14][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[14][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[14][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[14][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[14][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[14][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[14][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[14][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[14][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[14][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[14][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[14][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[14][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[14][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[14][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[14][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[14][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[14][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[14][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[14][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[14][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[14][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[14][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[14][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[14][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[14][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[14][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[14][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[14][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[14][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[14][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[14][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[14][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[14][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[14][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[14][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[14][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[14][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[14][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[14][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[14][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[15][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[15][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[15][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[15][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[15][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[15][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[15][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[15][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[15][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[15][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[15][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[15][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[15][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[15][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[15][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[15][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[15][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[15][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[15][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[15][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[15][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[15][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[15][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[15][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[15][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[15][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[15][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[15][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[15][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[15][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[15][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[15][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[15][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[15][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[15][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[15][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[15][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[15][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[15][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[15][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[15][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[16][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[16][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[16][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[16][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[16][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[16][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[16][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[16][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[16][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[16][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[16][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[16][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[16][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[16][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[16][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[16][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[16][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[16][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[16][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[16][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[16][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[16][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[16][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[16][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[16][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[16][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[16][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[16][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[16][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[16][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[16][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[16][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[16][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[16][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[16][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[16][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[16][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[16][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[16][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[16][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[16][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[17][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[17][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[17][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[17][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[17][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[17][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[17][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[17][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[17][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[17][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[17][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[17][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[17][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[17][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[17][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[17][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[17][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[17][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[17][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[17][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[17][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[17][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[17][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[17][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[17][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[17][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[17][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[17][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[17][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[17][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[17][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[17][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[17][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[17][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[17][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[17][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[17][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[17][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[17][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[17][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[17][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[18][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[18][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[18][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[18][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[18][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[18][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[18][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[18][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[18][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[18][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[18][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[18][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[18][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[18][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[18][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[18][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[18][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[18][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[18][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[18][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[18][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[18][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[18][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[18][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[18][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[18][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[18][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[18][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[18][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[18][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[18][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[18][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[18][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[18][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[18][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[18][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[18][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[18][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[18][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[18][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[18][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[19][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[19][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[19][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[19][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[19][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[19][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[19][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[19][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[19][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[19][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[19][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[19][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[19][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[19][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[19][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[19][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[19][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[19][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[19][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[19][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[19][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[19][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[19][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[19][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[19][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[19][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[19][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[19][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[19][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[19][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[19][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[19][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[19][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[19][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[19][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[19][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[19][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[19][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[19][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[19][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[19][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[20][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[20][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[20][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[20][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[20][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[20][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[20][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[20][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[20][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[20][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[20][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[20][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[20][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[20][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[20][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[20][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[20][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[20][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[20][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[20][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[20][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[20][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[20][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[20][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[20][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[20][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[20][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[20][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[20][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[20][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[20][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[20][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[20][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[20][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[20][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[20][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[20][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[20][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[20][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[20][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[20][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[21][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[21][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[21][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[21][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[21][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[21][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[21][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[21][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[21][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[21][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[21][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[21][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[21][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[21][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[21][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[21][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[21][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[21][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[21][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[21][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[21][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[21][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[21][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[21][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[21][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[21][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[21][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[21][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[21][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[21][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[21][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[21][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[21][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[21][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[21][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[21][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[21][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[21][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[21][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[21][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[21][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[22][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[22][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[22][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[22][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[22][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[22][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[22][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[22][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[22][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[22][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[22][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[22][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[22][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[22][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[22][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[22][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[22][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[22][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[22][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[22][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[22][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[22][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[22][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[22][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[22][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[22][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[22][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[22][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[22][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[22][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[22][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[22][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[22][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[22][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[22][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[22][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[22][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[22][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[22][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[22][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[22][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[23][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[23][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[23][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[23][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[23][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[23][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[23][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[23][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[23][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[23][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[23][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[23][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[23][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[23][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[23][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[23][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[23][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[23][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[23][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[23][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[23][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[23][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[23][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[23][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[23][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[23][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[23][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[23][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[23][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[23][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[23][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[23][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[23][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[23][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[23][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[23][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[23][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[23][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[23][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[23][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[23][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[24][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[24][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[24][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[24][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[24][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[24][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[24][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[24][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[24][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[24][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[24][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[24][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[24][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[24][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[24][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[24][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[24][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[24][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[24][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[24][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[24][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[24][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[24][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[24][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[24][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[24][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[24][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[24][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[24][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[24][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[24][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[24][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[24][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[24][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[24][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[24][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[24][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[24][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[24][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[24][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[24][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[25][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[25][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[25][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[25][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[25][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[25][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[25][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[25][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[25][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[25][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[25][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[25][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[25][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[25][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[25][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[25][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[25][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[25][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[25][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[25][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[25][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[25][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[25][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[25][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[25][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[25][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[25][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[25][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[25][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[25][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[25][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[25][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[25][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[25][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[25][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[25][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[25][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[25][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[25][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[25][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[25][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[26][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[26][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[26][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[26][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[26][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[26][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[26][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[26][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[26][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[26][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[26][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[26][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[26][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[26][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[26][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[26][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[26][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[26][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[26][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[26][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[26][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[26][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[26][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[26][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[26][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[26][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[26][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[26][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[26][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[26][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[26][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[26][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[26][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[26][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[26][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[26][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[26][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[26][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[26][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[26][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[26][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[27][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[27][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[27][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[27][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[27][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[27][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[27][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[27][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[27][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[27][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[27][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[27][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[27][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[27][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[27][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[27][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[27][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[27][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[27][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[27][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[27][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[27][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[27][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[27][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[27][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[27][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[27][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[27][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[27][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[27][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[27][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[27][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[27][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[27][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[27][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[27][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[27][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[27][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[27][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[27][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[27][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[28][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[28][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[28][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[28][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[28][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[28][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[28][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[28][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[28][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[28][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[28][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[28][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[28][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[28][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[28][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[28][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[28][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[28][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[28][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[28][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[28][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[28][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[28][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[28][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[28][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[28][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[28][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[28][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[28][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[28][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[28][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[28][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[28][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[28][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[28][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[28][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[28][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[28][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[28][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[28][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[28][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[29][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[29][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[29][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[29][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[29][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[29][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[29][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[29][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[29][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[29][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[29][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[29][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[29][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[29][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[29][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[29][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[29][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[29][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[29][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[29][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[29][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[29][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[29][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[29][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[29][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[29][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[29][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[29][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[29][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[29][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[29][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[29][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[29][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[29][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[29][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[29][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[29][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[29][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[29][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[29][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[29][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[30][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[30][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[30][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[30][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[30][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[30][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[30][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[30][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[30][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[30][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[30][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[30][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[30][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[30][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[30][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[30][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[30][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[30][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[30][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[30][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[30][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[30][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[30][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[30][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[30][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[30][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[30][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[30][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[30][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[30][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[30][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[30][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[30][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[30][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[30][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[30][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[30][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[30][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[30][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[30][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[30][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[31][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[31][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[31][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[31][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[31][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[31][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[31][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[31][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[31][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[31][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[31][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[31][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[31][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[31][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[31][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[31][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[31][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[31][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[31][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[31][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[31][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[31][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[31][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[31][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[31][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[31][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[31][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[31][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[31][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[31][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[31][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[31][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[31][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[31][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[31][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[31][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[31][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[31][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[31][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[31][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[31][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[32][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[32][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[32][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[32][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[32][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[32][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[32][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[32][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[32][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[32][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[32][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[32][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[32][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[32][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[32][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[32][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[32][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[32][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[32][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[32][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[32][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[32][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[32][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[32][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[32][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[32][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[32][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[32][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[32][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[32][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[32][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[32][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[32][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[32][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[32][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[32][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[32][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[32][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[32][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[32][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[32][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[33][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[33][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[33][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[33][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[33][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[33][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[33][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[33][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[33][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[33][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[33][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[33][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[33][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[33][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[33][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[33][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[33][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[33][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[33][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[33][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[33][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[33][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[33][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[33][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[33][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[33][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[33][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[33][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[33][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[33][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[33][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[33][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[33][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[33][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[33][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[33][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[33][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[33][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[33][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[33][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[33][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[34][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[34][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[34][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[34][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[34][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[34][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[34][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[34][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[34][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[34][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[34][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[34][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[34][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[34][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[34][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[34][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[34][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[34][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[34][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[34][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[34][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[34][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[34][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[34][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[34][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[34][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[34][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[34][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[34][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[34][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[34][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[34][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[34][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[34][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[34][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[34][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[34][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[34][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[34][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[34][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[34][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[35][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[35][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[35][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[35][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[35][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[35][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[35][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[35][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[35][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[35][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[35][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[35][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[35][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[35][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[35][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[35][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[35][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[35][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[35][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[35][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[35][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[35][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[35][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[35][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[35][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[35][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[35][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[35][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[35][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[35][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[35][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[35][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[35][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[35][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[35][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[35][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[35][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[35][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[35][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[35][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[35][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[36][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[36][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[36][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[36][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[36][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[36][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[36][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[36][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[36][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[36][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[36][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[36][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[36][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[36][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[36][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[36][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[36][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[36][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[36][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[36][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[36][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[36][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[36][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[36][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[36][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[36][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[36][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[36][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[36][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[36][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[36][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[36][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[36][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[36][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[36][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[36][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[36][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[36][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[36][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[36][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[36][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[37][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[37][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[37][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[37][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[37][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[37][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[37][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[37][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[37][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[37][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[37][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[37][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[37][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[37][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[37][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[37][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[37][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[37][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[37][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[37][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[37][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[37][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[37][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[37][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[37][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[37][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[37][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[37][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[37][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[37][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[37][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[37][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[37][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[37][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[37][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[37][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[37][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[37][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[37][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[37][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[37][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[38][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[38][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[38][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[38][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[38][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[38][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[38][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[38][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[38][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[38][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[38][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[38][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[38][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[38][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[38][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[38][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[38][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[38][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[38][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[38][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[38][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[38][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[38][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[38][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[38][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[38][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[38][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[38][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[38][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[38][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[38][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[38][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[38][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[38][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[38][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[38][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[38][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[38][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[38][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[38][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[38][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[39][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[39][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[39][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[39][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[39][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[39][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[39][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[39][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[39][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[39][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[39][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[39][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[39][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[39][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[39][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[39][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[39][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[39][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[39][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[39][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[39][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[39][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[39][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[39][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[39][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[39][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[39][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[39][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[39][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[39][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[39][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[39][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[39][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[39][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[39][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[39][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[39][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[39][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[39][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[39][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[39][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[40][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[40][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[40][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[40][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[40][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[40][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[40][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[40][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[40][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[40][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[40][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[40][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[40][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[40][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[40][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[40][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[40][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[40][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[40][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[40][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[40][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[40][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[40][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[40][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[40][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[40][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[40][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[40][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[40][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[40][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[40][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[40][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[40][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[40][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[40][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[40][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[40][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[40][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[40][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[40][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[40][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[41][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[41][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[41][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[41][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[41][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[41][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[41][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[41][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[41][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[41][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[41][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[41][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[41][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[41][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[41][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[41][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[41][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[41][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[41][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[41][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[41][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[41][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[41][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[41][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[41][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[41][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[41][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[41][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[41][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[41][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[41][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[41][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[41][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[41][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[41][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[41][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[41][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[41][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[41][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[41][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[41][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[42][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[42][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[42][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[42][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[42][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[42][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[42][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[42][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[42][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[42][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[42][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[42][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[42][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[42][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[42][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[42][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[42][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[42][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[42][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[42][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[42][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[42][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[42][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[42][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[42][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[42][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[42][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[42][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[42][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[42][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[42][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[42][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[42][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[42][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[42][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[42][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[42][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[42][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[42][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[42][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[42][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[43][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[43][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[43][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[43][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[43][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[43][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[43][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[43][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[43][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[43][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[43][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[43][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[43][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[43][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[43][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[43][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[43][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[43][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[43][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[43][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[43][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[43][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[43][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[43][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[43][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[43][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[43][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[43][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[43][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[43][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[43][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[43][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[43][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[43][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[43][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[43][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[43][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[43][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[43][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[43][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[43][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[44][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[44][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[44][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[44][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[44][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[44][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[44][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[44][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[44][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[44][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[44][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[44][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[44][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[44][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[44][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[44][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[44][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[44][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[44][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[44][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[44][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[44][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[44][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[44][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[44][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[44][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[44][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[44][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[44][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[44][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[44][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[44][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[44][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[44][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[44][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[44][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[44][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[44][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[44][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[44][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[44][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[45][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[45][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[45][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[45][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[45][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[45][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[45][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[45][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[45][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[45][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[45][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[45][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[45][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[45][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[45][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[45][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[45][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[45][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[45][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[45][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[45][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[45][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[45][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[45][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[45][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[45][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[45][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[45][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[45][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[45][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[45][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[45][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[45][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[45][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[45][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[45][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[45][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[45][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[45][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[45][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[45][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[46][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[46][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[46][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[46][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[46][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[46][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[46][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[46][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[46][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[46][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[46][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[46][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[46][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[46][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[46][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[46][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[46][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[46][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[46][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[46][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[46][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[46][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[46][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[46][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[46][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[46][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[46][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[46][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[46][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[46][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[46][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[46][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[46][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[46][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[46][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[46][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[46][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[46][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[46][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[46][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[46][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[47][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[47][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[47][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[47][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[47][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[47][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[47][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[47][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[47][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[47][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[47][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[47][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[47][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[47][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[47][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[47][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[47][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[47][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[47][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[47][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[47][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[47][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[47][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[47][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[47][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[47][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[47][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[47][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[47][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[47][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[47][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[47][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[47][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[47][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[47][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[47][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[47][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[47][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[47][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[47][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[47][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[48][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[48][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[48][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[48][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[48][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[48][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[48][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[48][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[48][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[48][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[48][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[48][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[48][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[48][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[48][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[48][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[48][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[48][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[48][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[48][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[48][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[48][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[48][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[48][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[48][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[48][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[48][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[48][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[48][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[48][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[48][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[48][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[48][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[48][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[48][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[48][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[48][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[48][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[48][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[48][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[48][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[49][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[49][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[49][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[49][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[49][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[49][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[49][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[49][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[49][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[49][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[49][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[49][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[49][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[49][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[49][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[49][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[49][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[49][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[49][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[49][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[49][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[49][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[49][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[49][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[49][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[49][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[49][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[49][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[49][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[49][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[49][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[49][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[49][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[49][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[49][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[49][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[49][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[49][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[49][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[49][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[49][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[50][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[50][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[50][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[50][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[50][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[50][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[50][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[50][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[50][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[50][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[50][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[50][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[50][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[50][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[50][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[50][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[50][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[50][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[50][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[50][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[50][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[50][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[50][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[50][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[50][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[50][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[50][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[50][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[50][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[50][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[50][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[50][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[50][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[50][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[50][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[50][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[50][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[50][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[50][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[50][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[50][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[51][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[51][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[51][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[51][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[51][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[51][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[51][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[51][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[51][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[51][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[51][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[51][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[51][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[51][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[51][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[51][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[51][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[51][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[51][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[51][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[51][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[51][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[51][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[51][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[51][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[51][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[51][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[51][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[51][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[51][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[51][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[51][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[51][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[51][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[51][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[51][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[51][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[51][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[51][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[51][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[51][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[52][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[52][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[52][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[52][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[52][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[52][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[52][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[52][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[52][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[52][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[52][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[52][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[52][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[52][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[52][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[52][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[52][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[52][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[52][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[52][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[52][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[52][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[52][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[52][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[52][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[52][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[52][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[52][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[52][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[52][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[52][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[52][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[52][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[52][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[52][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[52][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[52][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[52][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[52][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[52][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[52][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[53][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[53][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[53][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[53][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[53][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[53][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[53][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[53][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[53][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[53][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[53][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[53][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[53][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[53][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[53][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[53][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[53][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[53][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[53][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[53][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[53][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[53][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[53][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[53][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[53][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[53][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[53][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[53][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[53][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[53][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[53][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[53][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[53][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[53][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[53][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[53][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[53][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[53][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[53][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[53][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[53][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[54][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[54][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[54][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[54][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[54][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[54][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[54][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[54][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[54][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[54][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[54][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[54][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[54][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[54][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[54][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[54][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[54][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[54][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[54][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[54][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[54][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[54][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[54][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[54][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[54][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[54][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[54][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[54][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[54][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[54][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[54][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[54][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[54][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[54][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[54][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[54][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[54][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[54][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[54][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[54][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[54][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[55][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[55][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[55][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[55][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[55][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[55][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[55][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[55][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[55][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[55][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[55][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[55][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[55][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[55][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[55][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[55][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[55][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[55][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[55][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[55][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[55][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[55][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[55][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[55][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[55][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[55][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[55][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[55][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[55][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[55][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[55][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[55][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[55][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[55][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[55][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[55][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[55][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[55][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[55][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[55][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[55][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[56][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[56][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[56][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[56][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[56][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[56][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[56][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[56][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[56][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[56][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[56][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[56][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[56][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[56][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[56][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[56][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[56][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[56][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[56][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[56][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[56][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[56][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[56][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[56][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[56][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[56][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[56][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[56][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[56][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[56][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[56][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[56][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[56][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[56][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[56][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[56][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[56][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[56][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[56][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[56][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[56][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[57][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[57][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[57][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[57][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[57][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[57][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[57][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[57][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[57][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[57][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[57][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[57][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[57][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[57][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[57][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[57][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[57][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[57][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[57][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[57][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[57][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[57][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[57][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[57][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[57][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[57][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[57][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[57][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[57][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[57][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[57][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[57][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[57][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[57][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[57][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[57][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[57][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[57][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[57][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[57][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[57][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[58][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[58][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[58][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[58][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[58][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[58][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[58][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[58][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[58][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[58][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[58][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[58][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[58][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[58][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[58][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[58][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[58][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[58][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[58][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[58][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[58][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[58][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[58][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[58][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[58][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[58][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[58][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[58][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[58][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[58][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[58][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[58][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[58][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[58][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[58][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[58][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[58][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[58][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[58][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[58][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[58][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[59][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[59][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[59][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[59][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[59][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[59][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[59][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[59][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[59][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[59][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[59][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[59][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[59][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[59][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[59][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[59][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[59][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[59][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[59][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[59][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[59][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[59][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[59][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[59][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[59][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[59][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[59][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[59][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[59][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[59][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[59][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[59][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[59][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[59][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[59][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[59][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[59][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[59][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[59][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[59][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[59][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[60][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[60][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[60][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[60][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[60][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[60][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[60][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[60][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[60][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[60][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[60][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[60][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[60][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[60][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[60][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[60][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[60][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[60][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[60][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[60][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[60][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[60][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[60][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[60][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[60][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[60][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[60][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[60][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[60][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[60][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[60][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[60][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[60][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[60][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[60][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[60][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[60][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[60][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[60][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[60][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[60][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[61][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[61][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[61][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[61][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[61][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[61][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[61][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[61][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[61][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[61][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[61][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[61][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[61][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[61][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[61][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[61][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[61][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[61][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[61][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[61][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[61][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[61][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[61][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[61][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[61][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[61][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[61][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[61][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[61][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[61][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[61][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[61][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[61][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[61][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[61][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[61][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[61][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[61][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[61][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[61][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[61][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[62][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[62][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[62][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[62][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[62][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[62][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[62][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[62][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[62][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[62][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[62][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[62][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[62][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[62][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[62][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[62][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[62][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[62][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[62][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[62][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[62][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[62][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[62][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[62][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[62][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[62][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[62][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[62][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[62][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[62][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[62][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[62][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[62][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[62][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[62][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[62][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[62][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[62][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[62][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[62][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[62][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[63][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[63][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[63][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[63][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[63][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[63][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[63][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[63][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[63][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[63][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[63][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[63][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[63][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[63][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[63][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[63][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[63][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[63][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[63][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[63][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[63][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[63][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[63][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[63][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[63][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[63][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[63][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[63][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[63][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[63][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[63][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[63][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[63][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[63][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[63][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[63][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[63][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[63][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[63][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[63][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[63][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[64][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[64][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[64][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[64][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[64][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[64][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[64][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[64][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[64][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[64][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[64][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[64][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[64][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[64][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[64][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[64][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[64][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[64][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[64][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[64][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[64][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[64][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[64][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[64][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[64][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[64][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[64][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[64][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[64][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[64][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[64][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[64][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[64][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[64][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[64][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[64][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[64][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[64][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[64][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[64][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[64][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[65][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[65][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[65][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[65][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[65][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[65][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[65][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[65][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[65][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[65][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[65][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[65][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[65][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[65][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[65][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[65][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[65][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[65][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[65][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[65][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[65][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[65][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[65][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[65][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[65][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[65][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[65][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[65][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[65][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[65][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[65][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[65][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[65][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[65][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[65][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[65][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[65][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[65][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[65][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[65][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[65][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[66][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[66][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[66][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[66][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[66][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[66][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[66][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[66][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[66][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[66][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[66][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[66][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[66][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[66][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[66][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[66][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[66][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[66][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[66][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[66][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[66][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[66][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[66][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[66][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[66][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[66][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[66][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[66][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[66][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[66][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[66][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[66][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[66][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[66][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[66][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[66][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[66][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[66][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[66][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[66][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[66][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[67][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[67][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[67][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[67][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[67][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[67][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[67][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[67][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[67][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[67][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[67][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[67][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[67][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[67][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[67][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[67][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[67][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[67][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[67][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[67][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[67][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[67][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[67][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[67][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[67][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[67][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[67][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[67][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[67][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[67][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[67][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[67][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[67][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[67][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[67][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[67][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[67][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[67][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[67][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[67][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[67][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[68][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[68][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[68][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[68][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[68][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[68][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[68][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[68][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[68][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[68][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[68][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[68][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[68][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[68][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[68][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[68][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[68][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[68][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[68][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[68][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[68][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[68][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[68][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[68][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[68][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[68][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[68][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[68][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[68][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[68][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[68][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[68][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[68][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[68][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[68][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[68][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[68][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[68][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[68][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[68][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[68][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[69][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[69][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[69][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[69][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[69][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[69][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[69][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[69][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[69][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[69][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[69][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[69][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[69][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[69][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[69][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[69][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[69][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[69][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[69][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[69][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[69][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[69][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[69][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[69][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[69][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[69][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[69][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[69][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[69][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[69][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[69][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[69][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[69][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[69][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[69][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[69][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[69][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[69][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[69][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[69][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[69][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[70][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[70][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[70][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[70][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[70][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[70][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[70][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[70][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[70][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[70][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[70][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[70][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[70][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[70][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[70][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[70][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[70][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[70][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[70][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[70][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[70][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[70][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[70][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[70][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[70][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[70][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[70][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[70][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[70][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[70][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[70][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[70][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[70][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[70][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[70][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[70][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[70][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[70][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[70][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[70][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[70][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[71][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[71][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[71][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[71][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[71][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[71][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[71][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[71][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[71][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[71][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[71][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[71][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[71][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[71][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[71][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[71][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[71][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[71][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[71][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[71][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[71][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[71][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[71][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[71][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[71][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[71][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[71][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[71][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[71][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[71][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[71][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[71][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[71][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[71][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[71][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[71][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[71][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[71][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[71][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[71][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[71][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[72][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[72][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[72][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[72][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[72][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[72][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[72][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[72][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[72][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[72][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[72][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[72][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[72][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[72][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[72][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[72][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[72][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[72][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[72][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[72][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[72][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[72][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[72][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[72][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[72][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[72][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[72][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[72][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[72][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[72][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[72][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[72][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[72][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[72][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[72][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[72][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[72][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[72][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[72][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[72][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[72][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[73][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[73][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[73][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[73][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[73][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[73][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[73][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[73][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[73][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[73][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[73][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[73][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[73][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[73][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[73][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[73][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[73][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[73][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[73][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[73][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[73][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[73][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[73][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[73][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[73][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[73][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[73][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[73][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[73][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[73][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[73][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[73][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[73][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[73][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[73][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[73][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[73][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[73][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[73][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[73][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[73][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[74][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[74][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[74][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[74][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[74][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[74][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[74][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[74][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[74][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[74][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[74][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[74][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[74][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[74][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[74][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[74][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[74][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[74][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[74][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[74][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[74][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[74][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[74][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[74][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[74][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[74][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[74][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[74][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[74][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[74][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[74][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[74][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[74][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[74][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[74][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[74][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[74][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[74][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[74][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[74][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[74][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[75][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[75][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[75][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[75][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[75][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[75][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[75][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[75][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[75][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[75][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[75][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[75][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[75][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[75][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[75][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[75][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[75][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[75][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[75][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[75][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[75][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[75][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[75][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[75][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[75][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[75][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[75][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[75][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[75][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[75][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[75][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[75][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[75][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[75][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[75][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[75][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[75][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[75][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[75][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[75][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[75][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[76][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[76][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[76][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[76][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[76][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[76][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[76][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[76][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[76][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[76][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[76][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[76][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[76][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[76][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[76][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[76][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[76][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[76][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[76][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[76][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[76][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[76][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[76][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[76][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[76][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[76][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[76][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[76][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[76][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[76][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[76][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[76][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[76][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[76][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[76][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[76][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[76][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[76][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[76][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[76][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[76][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[77][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[77][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[77][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[77][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[77][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[77][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[77][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[77][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[77][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[77][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[77][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[77][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[77][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[77][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[77][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[77][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[77][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[77][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[77][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[77][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[77][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[77][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[77][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[77][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[77][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[77][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[77][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[77][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[77][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[77][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[77][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[77][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[77][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[77][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[77][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[77][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[77][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[77][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[77][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[77][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[77][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[78][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[78][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[78][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[78][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[78][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[78][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[78][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[78][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[78][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[78][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[78][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[78][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[78][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[78][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[78][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[78][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[78][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[78][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[78][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[78][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[78][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[78][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[78][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[78][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[78][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[78][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[78][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[78][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[78][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[78][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[78][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[78][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[78][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[78][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[78][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[78][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[78][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[78][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[78][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[78][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[78][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[79][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[79][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[79][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[79][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[79][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[79][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[79][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[79][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[79][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[79][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[79][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[79][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[79][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[79][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[79][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[79][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[79][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[79][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[79][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[79][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[79][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[79][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[79][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[79][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[79][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[79][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[79][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[79][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[79][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[79][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[79][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[79][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[79][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[79][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[79][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[79][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[79][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[79][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[79][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[79][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[79][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[80][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[80][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[80][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[80][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[80][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[80][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[80][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[80][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[80][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[80][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[80][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[80][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[80][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[80][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[80][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[80][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[80][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[80][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[80][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[80][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[80][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[80][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[80][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[80][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[80][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[80][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[80][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[80][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[80][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[80][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[80][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[80][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[80][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[80][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[80][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[80][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[80][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[80][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[80][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[80][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[80][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[81][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[81][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[81][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[81][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[81][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[81][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[81][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[81][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[81][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[81][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[81][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[81][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[81][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[81][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[81][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[81][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[81][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[81][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[81][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[81][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[81][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[81][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[81][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[81][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[81][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[81][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[81][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[81][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[81][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[81][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[81][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[81][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[81][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[81][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[81][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[81][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[81][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[81][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[81][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[81][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[81][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[82][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[82][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[82][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[82][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[82][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[82][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[82][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[82][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[82][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[82][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[82][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[82][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[82][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[82][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[82][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[82][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[82][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[82][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[82][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[82][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[82][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[82][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[82][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[82][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[82][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[82][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[82][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[82][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[82][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[82][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[82][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[82][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[82][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[82][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[82][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[82][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[82][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[82][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[82][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[82][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[82][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[83][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[83][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[83][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[83][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[83][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[83][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[83][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[83][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[83][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[83][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[83][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[83][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[83][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[83][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[83][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[83][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[83][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[83][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[83][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[83][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[83][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[83][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[83][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[83][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[83][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[83][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[83][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[83][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[83][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[83][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[83][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[83][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[83][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[83][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[83][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[83][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[83][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[83][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[83][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[83][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[83][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[84][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[84][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[84][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[84][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[84][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[84][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[84][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[84][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[84][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[84][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[84][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[84][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[84][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[84][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[84][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[84][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[84][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[84][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[84][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[84][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[84][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[84][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[84][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[84][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[84][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[84][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[84][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[84][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[84][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[84][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[84][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[84][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[84][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[84][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[84][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[84][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[84][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[84][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[84][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[84][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[84][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[85][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[85][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[85][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[85][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[85][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[85][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[85][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[85][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[85][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[85][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[85][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[85][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[85][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[85][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[85][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[85][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[85][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[85][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[85][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[85][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[85][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[85][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[85][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[85][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[85][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[85][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[85][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[85][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[85][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[85][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[85][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[85][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[85][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[85][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[85][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[85][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[85][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[85][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[85][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[85][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[85][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[86][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[86][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[86][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[86][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[86][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[86][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[86][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[86][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[86][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[86][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[86][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[86][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[86][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[86][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[86][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[86][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[86][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[86][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[86][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[86][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[86][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[86][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[86][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[86][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[86][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[86][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[86][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[86][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[86][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[86][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[86][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[86][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[86][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[86][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[86][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[86][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[86][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[86][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[86][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[86][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[86][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[87][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[87][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[87][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[87][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[87][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[87][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[87][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[87][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[87][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[87][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[87][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[87][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[87][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[87][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[87][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[87][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[87][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[87][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[87][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[87][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[87][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[87][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[87][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[87][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[87][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[87][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[87][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[87][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[87][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[87][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[87][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[87][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[87][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[87][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[87][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[87][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[87][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[87][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[87][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[87][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[87][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[88][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[88][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[88][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[88][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[88][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[88][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[88][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[88][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[88][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[88][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[88][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[88][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[88][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[88][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[88][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[88][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[88][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[88][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[88][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[88][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[88][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[88][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[88][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[88][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[88][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[88][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[88][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[88][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[88][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[88][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[88][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[88][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[88][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[88][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[88][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[88][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[88][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[88][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[88][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[88][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[88][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[89][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[89][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[89][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[89][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[89][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[89][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[89][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[89][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[89][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[89][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[89][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[89][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[89][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[89][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[89][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[89][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[89][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[89][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[89][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[89][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[89][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[89][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[89][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[89][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[89][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[89][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[89][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[89][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[89][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[89][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[89][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[89][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[89][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[89][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[89][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[89][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[89][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[89][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[89][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[89][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[89][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[90][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[90][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[90][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[90][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[90][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[90][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[90][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[90][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[90][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[90][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[90][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[90][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[90][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[90][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[90][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[90][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[90][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[90][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[90][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[90][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[90][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[90][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[90][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[90][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[90][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[90][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[90][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[90][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[90][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[90][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[90][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[90][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[90][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[90][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[90][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[90][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[90][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[90][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[90][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[90][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[90][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[91][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[91][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[91][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[91][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[91][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[91][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[91][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[91][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[91][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[91][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[91][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[91][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[91][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[91][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[91][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[91][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[91][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[91][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[91][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[91][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[91][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[91][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[91][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[91][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[91][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[91][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[91][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[91][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[91][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[91][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[91][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[91][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[91][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[91][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[91][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[91][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[91][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[91][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[91][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[91][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[91][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[92][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[92][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[92][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[92][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[92][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[92][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[92][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[92][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[92][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[92][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[92][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[92][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[92][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[92][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[92][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[92][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[92][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[92][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[92][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[92][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[92][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[92][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[92][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[92][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[92][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[92][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[92][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[92][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[92][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[92][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[92][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[92][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[92][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[92][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[92][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[92][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[92][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[92][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[92][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[92][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[92][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[93][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[93][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[93][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[93][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[93][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[93][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[93][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[93][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[93][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[93][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[93][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[93][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[93][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[93][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[93][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[93][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[93][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[93][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[93][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[93][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[93][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[93][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[93][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[93][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[93][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[93][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[93][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[93][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[93][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[93][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[93][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[93][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[93][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[93][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[93][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[93][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[93][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[93][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[93][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[93][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[93][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[94][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[94][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[94][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[94][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[94][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[94][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[94][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[94][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[94][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[94][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[94][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[94][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[94][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[94][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[94][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[94][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[94][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[94][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[94][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[94][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[94][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[94][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[94][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[94][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[94][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[94][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[94][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[94][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[94][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[94][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[94][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[94][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[94][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[94][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[94][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[94][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[94][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[94][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[94][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[94][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[94][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[95][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[95][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[95][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[95][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[95][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[95][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[95][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[95][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[95][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[95][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[95][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[95][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[95][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[95][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[95][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[95][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[95][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[95][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[95][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[95][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[95][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[95][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[95][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[95][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[95][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[95][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[95][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[95][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[95][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[95][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[95][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[95][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[95][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[95][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[95][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[95][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[95][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[95][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[95][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[95][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[95][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[96][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[96][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[96][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[96][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[96][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[96][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[96][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[96][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[96][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[96][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[96][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[96][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[96][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[96][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[96][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[96][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[96][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[96][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[96][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[96][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[96][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[96][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[96][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[96][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[96][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[96][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[96][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[96][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[96][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[96][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[96][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[96][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[96][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[96][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[96][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[96][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[96][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[96][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[96][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[96][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[96][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[97][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[97][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[97][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[97][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[97][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[97][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[97][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[97][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[97][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[97][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[97][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[97][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[97][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[97][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[97][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[97][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[97][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[97][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[97][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[97][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[97][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[97][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[97][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[97][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[97][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[97][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[97][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[97][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[97][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[97][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[97][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[97][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[97][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[97][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[97][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[97][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[97][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[97][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[97][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[97][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[97][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[98][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[98][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[98][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[98][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[98][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[98][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[98][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[98][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[98][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[98][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[98][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[98][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[98][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[98][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[98][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[98][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[98][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[98][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[98][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[98][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[98][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[98][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[98][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[98][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[98][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[98][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[98][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[98][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[98][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[98][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[98][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[98][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[98][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[98][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[98][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[98][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[98][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[98][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[98][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[98][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[98][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[99][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[99][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[99][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[99][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[99][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[99][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[99][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[99][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[99][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[99][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[99][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[99][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[99][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[99][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[99][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[99][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[99][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[99][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[99][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[99][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[99][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[99][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[99][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[99][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[99][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[99][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[99][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[99][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[99][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[99][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[99][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[99][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[99][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[99][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[99][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[99][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[99][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[99][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[99][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[99][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[99][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[100][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[100][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[100][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[100][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[100][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[100][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[100][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[100][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[100][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[100][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[100][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[100][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[100][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[100][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[100][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[100][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[100][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[100][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[100][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[100][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[100][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[100][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[100][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[100][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[100][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[100][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[100][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[100][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[100][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[100][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[100][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[100][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[100][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[100][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[100][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[100][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[100][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[100][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[100][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[100][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[100][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[101][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[101][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[101][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[101][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[101][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[101][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[101][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[101][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[101][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[101][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[101][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[101][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[101][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[101][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[101][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[101][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[101][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[101][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[101][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[101][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[101][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[101][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[101][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[101][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[101][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[101][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[101][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[101][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[101][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[101][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[101][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[101][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[101][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[101][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[101][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[101][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[101][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[101][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[101][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[101][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[101][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[102][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[102][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[102][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[102][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[102][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[102][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[102][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[102][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[102][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[102][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[102][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[102][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[102][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[102][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[102][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[102][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[102][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[102][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[102][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[102][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[102][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[102][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[102][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[102][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[102][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[102][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[102][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[102][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[102][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[102][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[102][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[102][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[102][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[102][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[102][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[102][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[102][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[102][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[102][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[102][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[102][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[103][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[103][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[103][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[103][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[103][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[103][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[103][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[103][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[103][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[103][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[103][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[103][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[103][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[103][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[103][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[103][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[103][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[103][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[103][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[103][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[103][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[103][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[103][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[103][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[103][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[103][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[103][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[103][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[103][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[103][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[103][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[103][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[103][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[103][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[103][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[103][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[103][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[103][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[103][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[103][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[103][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[104][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[104][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[104][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[104][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[104][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[104][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[104][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[104][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[104][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[104][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[104][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[104][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[104][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[104][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[104][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[104][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[104][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[104][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[104][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[104][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[104][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[104][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[104][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[104][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[104][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[104][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[104][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[104][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[104][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[104][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[104][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[104][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[104][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[104][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[104][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[104][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[104][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[104][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[104][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[104][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[104][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[105][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[105][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[105][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[105][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[105][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[105][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[105][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[105][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[105][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[105][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[105][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[105][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[105][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[105][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[105][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[105][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[105][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[105][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[105][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[105][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[105][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[105][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[105][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[105][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[105][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[105][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[105][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[105][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[105][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[105][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[105][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[105][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[105][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[105][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[105][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[105][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[105][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[105][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[105][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[105][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[105][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[106][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[106][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[106][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[106][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[106][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[106][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[106][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[106][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[106][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[106][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[106][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[106][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[106][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[106][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[106][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[106][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[106][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[106][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[106][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[106][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[106][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[106][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[106][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[106][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[106][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[106][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[106][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[106][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[106][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[106][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[106][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[106][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[106][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[106][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[106][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[106][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[106][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[106][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[106][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[106][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[106][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[107][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[107][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[107][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[107][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[107][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[107][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[107][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[107][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[107][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[107][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[107][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[107][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[107][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[107][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[107][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[107][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[107][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[107][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[107][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[107][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[107][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[107][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[107][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[107][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[107][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[107][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[107][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[107][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[107][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[107][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[107][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[107][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[107][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[107][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[107][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[107][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[107][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[107][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[107][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[107][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[107][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[108][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[108][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[108][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[108][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[108][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[108][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[108][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[108][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[108][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[108][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[108][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[108][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[108][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[108][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[108][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[108][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[108][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[108][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[108][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[108][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[108][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[108][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[108][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[108][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[108][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[108][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[108][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[108][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[108][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[108][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[108][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[108][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[108][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[108][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[108][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[108][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[108][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[108][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[108][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[108][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[108][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[109][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[109][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[109][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[109][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[109][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[109][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[109][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[109][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[109][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[109][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[109][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[109][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[109][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[109][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[109][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[109][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[109][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[109][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[109][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[109][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[109][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[109][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[109][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[109][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[109][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[109][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[109][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[109][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[109][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[109][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[109][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[109][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[109][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[109][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[109][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[109][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[109][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[109][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[109][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[109][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[109][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[110][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[110][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[110][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[110][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[110][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[110][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[110][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[110][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[110][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[110][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[110][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[110][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[110][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[110][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[110][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[110][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[110][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[110][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[110][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[110][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[110][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[110][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[110][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[110][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[110][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[110][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[110][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[110][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[110][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[110][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[110][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[110][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[110][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[110][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[110][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[110][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[110][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[110][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[110][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[110][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[110][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[111][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[111][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[111][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[111][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[111][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[111][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[111][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[111][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[111][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[111][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[111][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[111][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[111][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[111][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[111][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[111][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[111][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[111][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[111][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[111][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[111][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[111][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[111][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[111][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[111][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[111][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[111][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[111][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[111][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[111][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[111][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[111][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[111][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[111][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[111][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[111][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[111][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[111][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[111][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[111][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[111][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[112][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[112][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[112][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[112][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[112][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[112][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[112][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[112][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[112][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[112][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[112][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[112][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[112][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[112][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[112][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[112][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[112][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[112][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[112][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[112][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[112][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[112][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[112][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[112][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[112][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[112][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[112][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[112][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[112][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[112][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[112][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[112][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[112][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[112][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[112][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[112][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[112][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[112][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[112][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[112][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[112][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[113][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[113][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[113][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[113][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[113][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[113][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[113][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[113][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[113][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[113][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[113][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[113][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[113][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[113][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[113][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[113][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[113][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[113][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[113][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[113][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[113][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[113][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[113][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[113][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[113][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[113][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[113][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[113][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[113][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[113][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[113][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[113][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[113][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[113][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[113][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[113][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[113][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[113][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[113][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[113][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[113][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[114][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[114][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[114][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[114][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[114][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[114][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[114][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[114][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[114][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[114][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[114][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[114][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[114][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[114][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[114][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[114][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[114][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[114][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[114][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[114][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[114][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[114][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[114][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[114][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[114][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[114][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[114][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[114][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[114][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[114][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[114][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[114][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[114][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[114][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[114][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[114][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[114][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[114][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[114][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[114][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[114][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[115][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[115][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[115][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[115][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[115][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[115][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[115][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[115][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[115][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[115][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[115][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[115][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[115][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[115][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[115][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[115][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[115][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[115][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[115][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[115][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[115][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[115][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[115][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[115][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[115][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[115][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[115][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[115][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[115][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[115][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[115][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[115][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[115][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[115][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[115][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[115][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[115][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[115][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[115][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[115][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[115][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[116][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[116][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[116][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[116][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[116][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[116][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[116][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[116][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[116][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[116][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[116][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[116][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[116][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[116][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[116][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[116][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[116][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[116][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[116][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[116][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[116][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[116][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[116][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[116][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[116][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[116][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[116][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[116][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[116][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[116][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[116][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[116][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[116][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[116][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[116][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[116][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[116][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[116][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[116][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[116][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[116][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[117][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[117][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[117][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[117][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[117][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[117][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[117][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[117][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[117][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[117][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[117][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[117][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[117][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[117][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[117][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[117][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[117][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[117][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[117][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[117][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[117][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[117][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[117][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[117][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[117][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[117][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[117][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[117][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[117][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[117][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[117][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[117][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[117][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[117][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[117][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[117][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[117][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[117][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[117][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[117][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[117][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[118][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[118][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[118][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[118][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[118][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[118][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[118][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[118][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[118][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[118][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[118][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[118][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[118][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[118][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[118][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[118][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[118][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[118][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[118][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[118][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[118][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[118][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[118][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[118][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[118][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[118][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[118][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[118][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[118][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[118][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[118][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[118][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[118][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[118][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[118][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[118][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[118][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[118][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[118][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[118][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[118][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[119][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[119][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[119][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[119][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[119][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[119][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[119][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[119][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[119][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[119][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[119][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[119][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[119][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[119][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[119][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[119][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[119][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[119][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[119][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[119][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[119][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[119][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[119][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[119][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[119][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[119][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[119][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[119][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[119][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[119][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[119][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[119][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[119][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[119][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[119][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[119][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[119][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[119][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[119][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[119][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[119][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[120][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[120][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[120][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[120][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[120][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[120][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[120][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[120][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[120][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[120][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[120][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[120][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[120][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[120][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[120][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[120][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[120][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[120][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[120][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[120][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[120][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[120][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[120][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[120][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[120][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[120][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[120][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[120][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[120][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[120][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[120][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[120][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[120][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[120][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[120][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[120][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[120][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[120][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[120][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[120][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[120][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[121][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[121][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[121][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[121][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[121][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[121][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[121][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[121][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[121][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[121][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[121][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[121][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[121][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[121][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[121][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[121][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[121][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[121][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[121][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[121][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[121][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[121][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[121][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[121][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[121][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[121][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[121][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[121][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[121][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[121][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[121][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[121][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[121][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[121][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[121][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[121][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[121][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[121][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[121][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[121][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[121][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[122][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[122][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[122][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[122][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[122][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[122][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[122][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[122][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[122][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[122][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[122][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[122][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[122][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[122][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[122][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[122][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[122][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[122][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[122][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[122][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[122][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[122][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[122][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[122][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[122][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[122][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[122][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[122][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[122][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[122][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[122][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[122][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[122][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[122][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[122][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[122][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[122][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[122][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[122][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[122][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[122][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[123][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[123][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[123][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[123][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[123][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[123][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[123][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[123][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[123][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[123][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[123][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[123][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[123][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[123][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[123][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[123][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[123][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[123][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[123][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[123][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[123][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[123][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[123][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[123][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[123][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[123][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[123][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[123][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[123][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[123][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[123][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[123][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[123][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[123][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[123][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[123][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[123][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[123][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[123][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[123][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[123][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[124][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[124][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[124][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[124][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[124][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[124][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[124][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[124][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[124][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[124][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[124][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[124][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[124][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[124][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[124][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[124][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[124][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[124][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[124][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[124][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[124][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[124][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[124][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[124][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[124][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[124][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[124][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[124][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[124][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[124][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[124][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[124][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[124][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[124][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[124][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[124][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[124][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[124][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[124][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[124][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[124][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[125][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[125][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[125][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[125][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[125][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[125][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[125][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[125][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[125][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[125][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[125][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[125][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[125][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[125][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[125][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[125][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[125][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[125][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[125][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[125][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[125][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[125][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[125][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[125][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[125][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[125][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[125][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[125][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[125][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[125][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[125][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[125][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[125][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[125][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[125][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[125][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[125][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[125][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[125][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[125][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[125][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[126][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[126][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[126][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[126][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[126][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[126][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[126][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[126][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[126][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[126][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[126][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[126][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[126][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[126][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[126][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[126][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[126][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[126][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[126][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[126][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[126][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[126][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[126][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[126][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[126][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[126][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[126][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[126][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[126][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[126][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[126][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[126][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[126][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[126][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[126][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[126][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[126][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[126][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[126][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[126][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[126][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[127][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i11/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[127][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[127][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][0]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][0]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][0]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][0]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[127][0]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[127][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[127][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i11/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[127][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[127][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][1]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][1]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][1]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][1]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[127][1]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[127][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[127][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i11/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[127][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[127][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][2]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][2]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][2]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][2]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[127][2]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[127][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[127][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i11/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[127][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[127][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][3]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][3]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][3]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][3]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[127][3]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[127][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[127][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i11/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[127][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[127][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][4]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][4]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][4]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][4]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[127][4]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[127][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[127][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i11/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[127][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[127][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][5]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][5]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][5]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][5]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[127][5]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[127][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[127][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i11/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[127][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[127][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][6]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][6]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][6]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][6]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[127][6]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[127][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i11/fifo_inst/buff[127][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i11/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i11/fifo_inst/buff[127][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i11/fifo_inst/buff[127][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][7]~FF .CE_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][7]~FF .SR_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][7]~FF .D_POLARITY = 1'b1;
    defparam \i11/fifo_inst/buff[127][7]~FF .SR_SYNC = 1'b1;
    defparam \i11/fifo_inst/buff[127][7]~FF .SR_VALUE = 1'b0;
    defparam \i11/fifo_inst/buff[127][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \tx_dac_fsm_inst/i119  (.I0(n1417), .I1(n131), .I2(n1416), 
            .O(n131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/i119 .LUTMASK = 16'hacac;
    EFX_LUT4 \tx_dac_fsm_inst/dlatchrs_164/i1  (.I0(n1418), .I1(n132), .I2(n1416), 
            .O(n132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/dlatchrs_164/i1 .LUTMASK = 16'hacac;
    EFX_LUT4 \tx_dac_fsm_inst/dlatchrs_162/i2  (.I0(n1436), .I1(n150), .I2(n1411), 
            .O(n150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/dlatchrs_162/i2 .LUTMASK = 16'hacac;
    EFX_LUT4 \tx_dac_fsm_inst/dlatchrs_162/i3  (.I0(n1437), .I1(n151), .I2(n1411), 
            .O(n151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/dlatchrs_162/i3 .LUTMASK = 16'hacac;
    EFX_LUT4 \tx_dac_fsm_inst/dlatchrs_162/i4  (.I0(n1438), .I1(n152), .I2(n1411), 
            .O(n152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/dlatchrs_162/i4 .LUTMASK = 16'hacac;
    EFX_LUT4 \tx_dac_fsm_inst/dlatchrs_164/i2  (.I0(n1439), .I1(n153), .I2(n1416), 
            .O(n153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/dlatchrs_164/i2 .LUTMASK = 16'hacac;
    EFX_LUT4 LUT__2981 (.I0(\spi_slave_inst/bitcnt[4] ), .I1(\spi_slave_inst/bitcnt[3] ), 
            .O(n1703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__2981.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__2982 (.I0(n1703), .I1(rw_out), .I2(\spi_slave_inst/d_o[7] ), 
            .O(MISO)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__2982.LUTMASK = 16'h4040;
    EFX_ADD \led_inst/add_23/i2  (.I0(\led_inst/counter[1] ), .I1(\led_inst/counter[0] ), 
            .CI(1'b0), .O(n18), .CO(n19)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i2 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_129/i2  (.I0(\tx_dac_fsm_inst/zctr[1] ), 
            .I1(\tx_dac_fsm_inst/zctr[0] ), .CI(1'b0), .O(n135), .CO(n136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(197)
    defparam \tx_dac_fsm_inst/add_129/i2 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_129/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_136/i2  (.I0(\tx_dac_fsm_inst/dctr[1] ), 
            .I1(\tx_dac_fsm_inst/dctr[0] ), .CI(1'b0), .O(n138), .CO(n139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(208)
    defparam \tx_dac_fsm_inst/add_136/i2 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_136/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \fifo_inst/add_12/i2  (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[0] ), 
            .CI(1'b0), .O(n141), .CO(n142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(59)
    defparam \fifo_inst/add_12/i2 .I0_POLARITY = 1'b1;
    defparam \fifo_inst/add_12/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \fifo_inst/add_12/i8  (.I0(\fifo_inst/wr_index[7] ), .I1(1'b0), 
            .CI(n1071), .O(n1067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(59)
    defparam \fifo_inst/add_12/i8 .I0_POLARITY = 1'b1;
    defparam \fifo_inst/add_12/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \fifo_inst/add_12/i7  (.I0(\fifo_inst/wr_index[6] ), .I1(1'b0), 
            .CI(n1074), .O(n1070), .CO(n1071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(59)
    defparam \fifo_inst/add_12/i7 .I0_POLARITY = 1'b1;
    defparam \fifo_inst/add_12/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \fifo_inst/add_12/i6  (.I0(\fifo_inst/wr_index[5] ), .I1(1'b0), 
            .CI(n1078), .O(n1073), .CO(n1074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(59)
    defparam \fifo_inst/add_12/i6 .I0_POLARITY = 1'b1;
    defparam \fifo_inst/add_12/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \fifo_inst/add_12/i5  (.I0(\fifo_inst/wr_index[4] ), .I1(1'b0), 
            .CI(n1081), .O(n1077), .CO(n1078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(59)
    defparam \fifo_inst/add_12/i5 .I0_POLARITY = 1'b1;
    defparam \fifo_inst/add_12/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \fifo_inst/add_12/i4  (.I0(\fifo_inst/wr_index[3] ), .I1(1'b0), 
            .CI(n1084), .O(n1080), .CO(n1081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(59)
    defparam \fifo_inst/add_12/i4 .I0_POLARITY = 1'b1;
    defparam \fifo_inst/add_12/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \fifo_inst/add_12/i3  (.I0(\fifo_inst/wr_index[2] ), .I1(1'b0), 
            .CI(n142), .O(n1083), .CO(n1084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(59)
    defparam \fifo_inst/add_12/i3 .I0_POLARITY = 1'b1;
    defparam \fifo_inst/add_12/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_136/i6  (.I0(\tx_dac_fsm_inst/dctr[5] ), 
            .I1(1'b0), .CI(n1093), .O(n1090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(208)
    defparam \tx_dac_fsm_inst/add_136/i6 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_136/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_136/i5  (.I0(\tx_dac_fsm_inst/dctr[4] ), 
            .I1(1'b0), .CI(n1096), .O(n1092), .CO(n1093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(208)
    defparam \tx_dac_fsm_inst/add_136/i5 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_136/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_136/i4  (.I0(\tx_dac_fsm_inst/dctr[3] ), 
            .I1(1'b0), .CI(n2608), .O(n1095), .CO(n1096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(208)
    defparam \tx_dac_fsm_inst/add_136/i4 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_136/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_136/i3  (.I0(\tx_dac_fsm_inst/dctr[2] ), 
            .I1(1'b0), .CI(n139), .O(n1118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(208)
    defparam \tx_dac_fsm_inst/add_136/i3 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_136/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_129/i6  (.I0(\tx_dac_fsm_inst/zctr[5] ), 
            .I1(1'b0), .CI(n1127), .O(n1124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(197)
    defparam \tx_dac_fsm_inst/add_129/i6 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_129/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_129/i5  (.I0(\tx_dac_fsm_inst/zctr[4] ), 
            .I1(1'b0), .CI(n1131), .O(n1126), .CO(n1127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(197)
    defparam \tx_dac_fsm_inst/add_129/i5 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_129/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_129/i4  (.I0(\tx_dac_fsm_inst/zctr[3] ), 
            .I1(1'b0), .CI(n2609), .O(n1130), .CO(n1131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(197)
    defparam \tx_dac_fsm_inst/add_129/i4 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_129/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_129/i3  (.I0(\tx_dac_fsm_inst/zctr[2] ), 
            .I1(1'b0), .CI(n136), .O(n1133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(197)
    defparam \tx_dac_fsm_inst/add_129/i3 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_129/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/sub_20/add_2/i5  (.I0(\tx_dac_fsm_inst/sym_ctr[4] ), 
            .I1(1'b0), .CI(n2610), .O(n1139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(97)
    defparam \tx_dac_fsm_inst/sub_20/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sub_20/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/sub_20/add_2/i4  (.I0(\tx_dac_fsm_inst/sym_ctr[3] ), 
            .I1(1'b1), .CI(n2611), .O(n1141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(97)
    defparam \tx_dac_fsm_inst/sub_20/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sub_20/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_18/i5  (.I0(\tx_dac_fsm_inst/sym_ctr[4] ), 
            .I1(1'b0), .CI(n1154), .O(n1150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(95)
    defparam \tx_dac_fsm_inst/add_18/i5 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_18/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_18/i4  (.I0(\tx_dac_fsm_inst/sym_ctr[3] ), 
            .I1(1'b0), .CI(n1157), .O(n1153), .CO(n1154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(95)
    defparam \tx_dac_fsm_inst/add_18/i4 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_18/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_18/i3  (.I0(\tx_dac_fsm_inst/sym_ctr[2] ), 
            .I1(1'b0), .CI(n1160), .O(n1156), .CO(n1157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(95)
    defparam \tx_dac_fsm_inst/add_18/i3 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_18/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_18/i2  (.I0(\tx_dac_fsm_inst/sym_ctr[1] ), 
            .I1(1'b1), .CI(n2612), .O(n1159), .CO(n1160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(95)
    defparam \tx_dac_fsm_inst/add_18/i2 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_18/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i24  (.I0(\led_inst/counter[23] ), .I1(1'b0), 
            .CI(n1170), .O(n1167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i24 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i23  (.I0(\led_inst/counter[22] ), .I1(1'b0), 
            .CI(n1173), .O(n1169), .CO(n1170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i23 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i22  (.I0(\led_inst/counter[21] ), .I1(1'b0), 
            .CI(n1177), .O(n1172), .CO(n1173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i22 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i21  (.I0(\led_inst/counter[20] ), .I1(1'b0), 
            .CI(n1180), .O(n1176), .CO(n1177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i21 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i20  (.I0(\led_inst/counter[19] ), .I1(1'b0), 
            .CI(n1183), .O(n1179), .CO(n1180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i20 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i19  (.I0(\led_inst/counter[18] ), .I1(1'b0), 
            .CI(n1187), .O(n1182), .CO(n1183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i19 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i18  (.I0(\led_inst/counter[17] ), .I1(1'b0), 
            .CI(n1190), .O(n1186), .CO(n1187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i18 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i17  (.I0(\led_inst/counter[16] ), .I1(1'b0), 
            .CI(n1193), .O(n1189), .CO(n1190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i17 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i16  (.I0(\led_inst/counter[15] ), .I1(1'b0), 
            .CI(n1197), .O(n1192), .CO(n1193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i16 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i15  (.I0(\led_inst/counter[14] ), .I1(1'b0), 
            .CI(n1206), .O(n1196), .CO(n1197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i15 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i14  (.I0(\led_inst/counter[13] ), .I1(1'b0), 
            .CI(n1210), .O(n1205), .CO(n1206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i14 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i13  (.I0(\led_inst/counter[12] ), .I1(1'b0), 
            .CI(n1220), .O(n1209), .CO(n1210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i13 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i12  (.I0(\led_inst/counter[11] ), .I1(1'b0), 
            .CI(n1225), .O(n1219), .CO(n1220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i12 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i11  (.I0(\led_inst/counter[10] ), .I1(1'b0), 
            .CI(n1229), .O(n1224), .CO(n1225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i11 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i10  (.I0(\led_inst/counter[9] ), .I1(1'b0), 
            .CI(n1233), .O(n1228), .CO(n1229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i10 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i9  (.I0(\led_inst/counter[8] ), .I1(1'b0), 
            .CI(n1238), .O(n1232), .CO(n1233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i9 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i8  (.I0(\led_inst/counter[7] ), .I1(1'b0), 
            .CI(n1242), .O(n1237), .CO(n1238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i8 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i7  (.I0(\led_inst/counter[6] ), .I1(1'b0), 
            .CI(n1248), .O(n1241), .CO(n1242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i7 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i6  (.I0(\led_inst/counter[5] ), .I1(1'b0), 
            .CI(n1252), .O(n1247), .CO(n1248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i6 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i5  (.I0(\led_inst/counter[4] ), .I1(1'b0), 
            .CI(n1255), .O(n1251), .CO(n1252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i5 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i4  (.I0(\led_inst/counter[3] ), .I1(1'b0), 
            .CI(n1259), .O(n1254), .CO(n1255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i4 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i3  (.I0(\led_inst/counter[2] ), .I1(1'b0), 
            .CI(n19), .O(n1258), .CO(n1259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i3 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \spi_slave_inst/add_29/i5  (.I0(\spi_slave_inst/bitcnt[4] ), .I1(1'b0), 
            .CI(n1268), .O(n1264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/add_29/i5 .I0_POLARITY = 1'b1;
    defparam \spi_slave_inst/add_29/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \spi_slave_inst/add_29/i4  (.I0(\spi_slave_inst/bitcnt[3] ), .I1(1'b0), 
            .CI(n1274), .O(n1267), .CO(n1268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/add_29/i4 .I0_POLARITY = 1'b1;
    defparam \spi_slave_inst/add_29/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \spi_slave_inst/add_29/i3  (.I0(\spi_slave_inst/bitcnt[2] ), .I1(1'b0), 
            .CI(n1278), .O(n1273), .CO(n1274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/add_29/i3 .I0_POLARITY = 1'b1;
    defparam \spi_slave_inst/add_29/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \spi_slave_inst/add_29/i2  (.I0(\spi_slave_inst/bitcnt[1] ), .I1(\spi_slave_inst/bitcnt[0] ), 
            .CI(1'b0), .O(n1277), .CO(n1278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/add_29/i2 .I0_POLARITY = 1'b1;
    defparam \spi_slave_inst/add_29/i2 .I1_POLARITY = 1'b1;
    EFX_LUT4 LUT__2983 (.I0(\gpo_inst/gp_config_reg[6] ), .I1(\gpo_inst/gp_config_reg[7] ), 
            .O(gpo_pins[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2983.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2984 (.I0(\gpo_inst/gp_config_reg[5] ), .I1(\gpo_inst/gp_config_reg[7] ), 
            .O(gpo_pins[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2984.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2985 (.I0(\gpo_inst/gp_config_reg[4] ), .I1(\gpo_inst/gp_config_reg[7] ), 
            .O(gpo_pins[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2985.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2986 (.I0(\gpo_inst/gp_config_reg[3] ), .I1(\gpo_inst/gp_config_reg[7] ), 
            .O(gpo_pins[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2986.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2987 (.I0(\gpo_inst/gp_config_reg[2] ), .I1(\gpo_inst/gp_config_reg[7] ), 
            .O(gpo_pins[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2987.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2988 (.I0(\gpo_inst/gp_config_reg[1] ), .I1(\gpo_inst/gp_config_reg[7] ), 
            .O(gpo_pins[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2988.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2989 (.I0(\gpo_inst/gp_config_reg[0] ), .I1(\gpo_inst/gp_config_reg[7] ), 
            .O(gpo_pins[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2989.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2990 (.I0(\tx_dac_fsm_inst/dac_config_reg[0] ), .I1(n153), 
            .O(lvds_tx_inst1_DATA[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2990.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2991 (.I0(n132), .I1(\tx_dac_fsm_inst/dac_config_reg[0] ), 
            .O(lvds_tx_inst1_DATA[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2991.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2992 (.I0(\spi_slave_inst/sync_ss[1] ), .I1(\spi_slave_inst/sync_ss[2] ), 
            .O(n1704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2992.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2993 (.I0(n1704), .I1(\reg_addr[2] ), .O(\spi_slave_inst/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2993.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2994 (.I0(\spi_slave_inst/bitcnt[2] ), .I1(\spi_slave_inst/bitcnt[1] ), 
            .I2(\spi_slave_inst/bitcnt[0] ), .O(n1705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__2994.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__2995 (.I0(\spi_slave_inst/sync_sclk[2] ), .I1(\spi_slave_inst/sync_ss[1] ), 
            .I2(\spi_slave_inst/sync_sclk[1] ), .O(n1706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__2995.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__2996 (.I0(n1705), .I1(n1706), .I2(n1703), .I3(n1704), 
            .O(ceg_net5)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__2996.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__2997 (.I0(n1704), .I1(\reg_addr[1] ), .O(\spi_slave_inst/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2997.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2998 (.I0(n1704), .I1(n1273), .O(\spi_slave_inst/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2998.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2999 (.I0(n1704), .I1(n1706), .O(ceg_net37)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__2999.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3000 (.I0(n1704), .I1(n1277), .O(\spi_slave_inst/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3000.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3001 (.I0(n1704), .I1(\reg_addr[0] ), .O(\spi_slave_inst/n97 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3001.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3002 (.I0(\reg_addr[0] ), .I1(\reg_addr[3] ), .I2(\reg_addr[1] ), 
            .I3(\reg_addr[2] ), .O(n1707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__3002.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__3003 (.I0(n1707), .I1(rw_out), .I2(addr_dv), .O(tx_en)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3003.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3004 (.I0(n1704), .I1(\spi_slave_inst/bitcnt[0] ), .O(\spi_slave_inst/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3004.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3005 (.I0(\spi_slave_inst/sync_ss[1] ), .I1(\spi_slave_inst/sync_ss[2] ), 
            .O(\spi_slave_inst/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3005.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3006 (.I0(\spi_slave_inst/n68 ), .I1(\spi_slave_inst/sync_mosi[1] ), 
            .O(\spi_slave_inst/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3006.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3007 (.I0(n1706), .I1(n1703), .I2(n1705), .I3(\spi_slave_inst/n68 ), 
            .O(ceg_net20)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__3007.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__3008 (.I0(n1704), .I1(\spi_slave_inst/sync_mosi[1] ), 
            .O(\spi_slave_inst/n98 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3008.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3009 (.I0(\reg_addr[2] ), .I1(\reg_addr[1] ), .I2(\reg_addr[3] ), 
            .O(n1708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3009.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3010 (.I0(n1708), .I1(rw_out), .I2(\reg_addr[0] ), .I3(addr_dv), 
            .O(n1709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3010.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3011 (.I0(\reg_addr[0] ), .I1(rw_out), .I2(n1708), .I3(addr_dv), 
            .O(tx_en_fifo)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__3011.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__3012 (.I0(\reg_addr[2] ), .I1(\reg_addr[1] ), .O(n1710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3012.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3013 (.I0(\tx_dac_fsm_inst/dac_config_reg[0] ), .I1(\data_from_led[0] ), 
            .I2(\reg_addr[0] ), .O(n1711)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3013.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3014 (.I0(n1711), .I1(n1710), .I2(rw_out), .I3(addr_dv), 
            .O(n1712)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__3014.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__3015 (.I0(tx_en_fifo), .I1(\fifo_inst/buff_head[0] ), 
            .I2(n1712), .O(n1713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__3015.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__3016 (.I0(n1709), .I1(\fifo_inst/length[0] ), .I2(n1713), 
            .O(n1714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3016.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3017 (.I0(n1714), .I1(\spi_slave_inst/sync_tx_en[1] ), 
            .I2(\spi_slave_inst/sync_tx_en[0] ), .O(\spi_slave_inst/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3017.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3018 (.I0(\spi_slave_inst/sync_tx_en[1] ), .I1(\spi_slave_inst/sync_tx_en[0] ), 
            .I2(n1706), .I3(tx_en), .O(ceg_net77)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__3018.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__3019 (.I0(rw_out), .I1(n1703), .I2(n1706), .I3(n1704), 
            .O(ceg_net98)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__3019.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__3020 (.I0(\spi_slave_inst/bitcnt[2] ), .I1(\spi_slave_inst/bitcnt[1] ), 
            .I2(\spi_slave_inst/bitcnt[0] ), .O(n1715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3020.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3021 (.I0(\spi_slave_inst/n68 ), .I1(n1715), .I2(n1703), 
            .O(ceg_net31)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3021.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3022 (.I0(\spi_slave_inst/bitcnt[4] ), .I1(\spi_slave_inst/sync_sclk[2] ), 
            .I2(\spi_slave_inst/sync_sclk[1] ), .I3(\spi_slave_inst/bitcnt[3] ), 
            .O(n1716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__3022.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__3023 (.I0(rw_out), .I1(n1715), .I2(n1716), .I3(\spi_slave_inst/n68 ), 
            .O(ceg_net34)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__3023.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__3024 (.I0(n1704), .I1(n1264), .O(\spi_slave_inst/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3024.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3025 (.I0(n1704), .I1(n1267), .O(\spi_slave_inst/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3025.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3026 (.I0(\reg_addr[0] ), .I1(rw_out), .I2(n1710), .I3(addr_dv), 
            .O(n1717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__3026.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__3027 (.I0(tx_en_fifo), .I1(n1717), .I2(\spi_slave_inst/sync_tx_en[1] ), 
            .I3(\spi_slave_inst/sync_tx_en[0] ), .O(n1718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__3027.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__3028 (.I0(n1718), .I1(\fifo_inst/buff_head[1] ), .I2(\fifo_inst/length[1] ), 
            .I3(n1709), .O(n1719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3028.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3029 (.I0(n1718), .I1(tx_en), .I2(n1706), .O(n1720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3029.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3030 (.I0(n1720), .I1(\spi_slave_inst/d_o[0] ), .I2(n1718), 
            .I3(\data_from_led[1] ), .O(n1721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3030.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3031 (.I0(n1717), .I1(\spi_slave_inst/sync_tx_en[1] ), 
            .I2(\spi_slave_inst/sync_tx_en[0] ), .O(n1722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3031.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3032 (.I0(n1721), .I1(n1719), .I2(n1722), .O(\spi_slave_inst/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3032.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3033 (.I0(n1718), .I1(\fifo_inst/buff_head[2] ), .I2(\fifo_inst/length[2] ), 
            .I3(n1709), .O(n1723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3033.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3034 (.I0(n1720), .I1(\spi_slave_inst/d_o[1] ), .I2(n1718), 
            .I3(\data_from_led[2] ), .O(n1724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3034.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3035 (.I0(n1724), .I1(n1723), .I2(n1722), .O(\spi_slave_inst/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3035.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3036 (.I0(n1718), .I1(\fifo_inst/buff_head[3] ), .I2(\fifo_inst/length[3] ), 
            .I3(n1709), .O(n1725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3036.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3037 (.I0(n1720), .I1(\spi_slave_inst/d_o[2] ), .I2(n1718), 
            .I3(\data_from_led[3] ), .O(n1726)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3037.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3038 (.I0(n1726), .I1(n1725), .I2(n1722), .O(\spi_slave_inst/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3038.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3039 (.I0(n1718), .I1(\fifo_inst/buff_head[4] ), .I2(\fifo_inst/length[4] ), 
            .I3(n1709), .O(n1727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3039.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3040 (.I0(n1720), .I1(\spi_slave_inst/d_o[3] ), .I2(n1718), 
            .I3(\data_from_led[4] ), .O(n1728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3040.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3041 (.I0(n1728), .I1(n1727), .I2(n1722), .O(\spi_slave_inst/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3041.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3042 (.I0(n1709), .I1(\fifo_inst/length[5] ), .I2(tx_en_fifo), 
            .I3(\fifo_inst/buff_head[5] ), .O(n1729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3042.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3043 (.I0(n1720), .I1(\spi_slave_inst/d_o[4] ), .I2(n1718), 
            .I3(\data_from_led[5] ), .O(n1730)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3043.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3044 (.I0(n1730), .I1(n1729), .I2(n1722), .O(\spi_slave_inst/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3044.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3045 (.I0(n1709), .I1(\fifo_inst/length[6] ), .I2(tx_en_fifo), 
            .I3(\fifo_inst/buff_head[6] ), .O(n1731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3045.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3046 (.I0(n1720), .I1(\spi_slave_inst/d_o[5] ), .I2(n1718), 
            .I3(\data_from_led[6] ), .O(n1732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3046.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3047 (.I0(n1732), .I1(n1731), .I2(n1722), .O(\spi_slave_inst/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3047.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3048 (.I0(n1709), .I1(\fifo_inst/length[7] ), .I2(tx_en_fifo), 
            .I3(\fifo_inst/buff_head[7] ), .O(n1733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3048.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3049 (.I0(n1720), .I1(\spi_slave_inst/d_o[6] ), .I2(n1718), 
            .I3(\data_from_led[7] ), .O(n1734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__3049.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__3050 (.I0(n1734), .I1(n1733), .I2(n1722), .O(\spi_slave_inst/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3050.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3051 (.I0(n1704), .I1(\rx_d[0] ), .O(\spi_slave_inst/n173 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3051.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3052 (.I0(n1704), .I1(\rx_d[1] ), .O(\spi_slave_inst/n172 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3052.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3053 (.I0(n1704), .I1(\rx_d[2] ), .O(\spi_slave_inst/n171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3053.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3054 (.I0(n1704), .I1(\rx_d[3] ), .O(\spi_slave_inst/n170 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3054.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3055 (.I0(n1704), .I1(\rx_d[4] ), .O(\spi_slave_inst/n169 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3055.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3056 (.I0(n1704), .I1(\rx_d[5] ), .O(\spi_slave_inst/n168 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3056.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3057 (.I0(n1704), .I1(\rx_d[6] ), .O(\spi_slave_inst/n167 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3057.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3058 (.I0(n1717), .I1(\led_inst/ctr_cfg_reg[7] ), .O(\led_inst/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3058.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3059 (.I0(n1717), .I1(\led_inst/ctr_cfg_reg[6] ), .O(\led_inst/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3059.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3060 (.I0(n1717), .I1(\led_inst/ctr_cfg_reg[5] ), .O(\led_inst/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3060.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3061 (.I0(n1717), .I1(\led_inst/ctr_cfg_reg[4] ), .O(\led_inst/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3061.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3062 (.I0(n1717), .I1(\led_inst/ctr_cfg_reg[3] ), .O(\led_inst/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3062.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3063 (.I0(n1717), .I1(\led_inst/ctr_cfg_reg[0] ), .O(\led_inst/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3063.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3064 (.I0(n1717), .I1(\led_inst/ctr_cfg_reg[2] ), .O(\led_inst/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3064.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3065 (.I0(n1717), .I1(\led_inst/ctr_cfg_reg[1] ), .O(\led_inst/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3065.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3066 (.I0(\led_inst/counter[17] ), .I1(\led_inst/counter[16] ), 
            .I2(\led_inst/ctr_cfg_reg[1] ), .I3(\led_inst/ctr_cfg_reg[0] ), 
            .O(n1735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__3066.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__3067 (.I0(n1735), .I1(\led_inst/ctr_cfg_reg[2] ), .I2(\led_inst/counter[18] ), 
            .O(n1736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__3067.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__3068 (.I0(\led_inst/ctr_cfg_reg[4] ), .I1(\led_inst/counter[20] ), 
            .O(n1737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3068.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3069 (.I0(n1736), .I1(\led_inst/counter[19] ), .I2(\led_inst/ctr_cfg_reg[3] ), 
            .I3(n1737), .O(n1738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0071 */ ;
    defparam LUT__3069.LUTMASK = 16'h0071;
    EFX_LUT4 LUT__3070 (.I0(\led_inst/counter[20] ), .I1(\led_inst/ctr_cfg_reg[4] ), 
            .O(n1739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3070.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3071 (.I0(\led_inst/counter[21] ), .I1(\led_inst/ctr_cfg_reg[5] ), 
            .I2(n1738), .I3(n1739), .O(n1740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hddd4 */ ;
    defparam LUT__3071.LUTMASK = 16'hddd4;
    EFX_LUT4 LUT__3072 (.I0(\led_inst/counter[22] ), .I1(\led_inst/ctr_cfg_reg[6] ), 
            .O(n1741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3072.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3073 (.I0(\led_inst/ctr_cfg_reg[6] ), .I1(\led_inst/counter[22] ), 
            .I2(\led_inst/ctr_cfg_reg[7] ), .I3(\led_inst/counter[23] ), 
            .O(n1742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__3073.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__3074 (.I0(\led_inst/counter[23] ), .I1(\led_inst/ctr_cfg_reg[7] ), 
            .O(n1743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3074.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3075 (.I0(n1741), .I1(n1740), .I2(n1742), .I3(n1743), 
            .O(\led_inst/LessThan_21/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__3075.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__3076 (.I0(\led_inst/LessThan_21/n48 ), .I1(\led_inst/counter[0] ), 
            .O(\led_inst/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3076.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3077 (.I0(rw_out), .I1(addr_dv), .I2(rxdv), .O(n1744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3077.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3078 (.I0(\reg_addr[0] ), .I1(n1744), .I2(n1710), .O(rx_en_led)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3078.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3079 (.I0(rx_en_led), .I1(\rx_d[0] ), .O(\data_to_led[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3079.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3080 (.I0(\led_inst/LessThan_21/n48 ), .I1(n18), .O(\led_inst/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3080.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3081 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1258), .O(\led_inst/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3081.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3082 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1254), .O(\led_inst/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3082.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3083 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1251), .O(\led_inst/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3083.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3084 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1247), .O(\led_inst/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3084.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3085 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1241), .O(\led_inst/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3085.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3086 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1237), .O(\led_inst/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3086.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3087 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1232), .O(\led_inst/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3087.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3088 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1228), .O(\led_inst/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3088.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3089 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1224), .O(\led_inst/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3089.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3090 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1219), .O(\led_inst/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3090.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3091 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1209), .O(\led_inst/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3091.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3092 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1205), .O(\led_inst/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3092.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3093 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1196), .O(\led_inst/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3093.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3094 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1192), .O(\led_inst/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3094.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3095 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1189), .O(\led_inst/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3095.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3096 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1186), .O(\led_inst/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3096.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3097 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1182), .O(\led_inst/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3097.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3098 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1179), .O(\led_inst/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3098.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3099 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1176), .O(\led_inst/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3099.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3100 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1172), .O(\led_inst/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3100.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3101 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1169), .O(\led_inst/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3101.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3102 (.I0(\led_inst/LessThan_21/n48 ), .I1(n1167), .O(\led_inst/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3102.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3103 (.I0(rx_en_led), .I1(\rx_d[1] ), .O(\data_to_led[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3103.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3104 (.I0(rx_en_led), .I1(\rx_d[2] ), .O(\data_to_led[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3104.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3105 (.I0(rx_en_led), .I1(\rx_d[3] ), .O(\data_to_led[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3105.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3106 (.I0(rx_en_led), .I1(\rx_d[4] ), .O(\data_to_led[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3106.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3107 (.I0(rx_en_led), .I1(\rx_d[5] ), .O(\data_to_led[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3107.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3108 (.I0(rx_en_led), .I1(\rx_d[6] ), .O(\data_to_led[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3108.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3109 (.I0(rx_en_led), .I1(\rx_d[7] ), .O(\data_to_led[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3109.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3110 (.I0(\reg_addr[2] ), .I1(\reg_addr[1] ), .I2(\reg_addr[0] ), 
            .I3(n1744), .O(rx_en_gpo)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3110.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3111 (.I0(rx_en_gpo), .I1(\reg_addr[3] ), .O(rx_en_fifo)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3111.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3112 (.I0(rx_en_fifo), .I1(\rx_d[5] ), .O(\data_to_fifo[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3112.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3113 (.I0(\fifo_inst/sync_wr[1] ), .I1(\fifo_inst/sync_wr[0] ), 
            .O(n1745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3113.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3114 (.I0(\fifo_inst/wr_index[0] ), .I1(\fifo_inst/wr_index[7] ), 
            .I2(n1745), .O(n1746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3114.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3115 (.I0(\fifo_inst/wr_index[5] ), .I1(\fifo_inst/wr_index[6] ), 
            .I2(n1746), .O(n1747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3115.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3116 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[3] ), 
            .I2(\fifo_inst/wr_index[4] ), .I3(\fifo_inst/wr_index[2] ), 
            .O(n1748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3116.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3117 (.I0(n1747), .I1(n1748), .O(\i11/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3117.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3118 (.I0(rx_en_gpo), .I1(\rx_d[0] ), .O(\data_to_gpo[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3118.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3119 (.I0(rx_en_fifo), .I1(\rx_d[4] ), .O(\data_to_fifo[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3119.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3120 (.I0(rx_en_gpo), .I1(\rx_d[1] ), .O(\data_to_gpo[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3120.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3121 (.I0(rx_en_gpo), .I1(\rx_d[2] ), .O(\data_to_gpo[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3121.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3122 (.I0(rx_en_gpo), .I1(\rx_d[3] ), .O(\data_to_gpo[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3122.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3123 (.I0(rx_en_gpo), .I1(\rx_d[4] ), .O(\data_to_gpo[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3123.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3124 (.I0(rx_en_gpo), .I1(\rx_d[5] ), .O(\data_to_gpo[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3124.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3125 (.I0(rx_en_gpo), .I1(\rx_d[6] ), .O(\data_to_gpo[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3125.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3126 (.I0(rx_en_gpo), .I1(\rx_d[7] ), .O(\data_to_gpo[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3126.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3127 (.I0(rx_en_fifo), .I1(\rx_d[0] ), .O(\data_to_fifo[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3127.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3128 (.I0(\fifo_inst/wr_index[2] ), .I1(\fifo_inst/wr_index[3] ), 
            .I2(\fifo_inst/wr_index[4] ), .I3(\fifo_inst/wr_index[1] ), 
            .O(n1749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3128.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3129 (.I0(n1747), .I1(n1749), .O(\i11/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3129.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3130 (.I0(rx_en_fifo), .I1(\rx_d[3] ), .O(\data_to_fifo[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3130.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3131 (.I0(rx_en_fifo), .I1(\rx_d[7] ), .O(\data_to_fifo[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3131.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3132 (.I0(\fifo_inst/wr_index[7] ), .I1(\fifo_inst/wr_index[0] ), 
            .I2(n1745), .O(n1750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3132.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3133 (.I0(\fifo_inst/wr_index[5] ), .I1(\fifo_inst/wr_index[6] ), 
            .I2(n1750), .O(n1751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3133.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3134 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[2] ), 
            .I2(\fifo_inst/wr_index[3] ), .I3(\fifo_inst/wr_index[4] ), 
            .O(n1752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3134.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3135 (.I0(n1751), .I1(n1752), .O(\i11/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3135.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3136 (.I0(rx_en_fifo), .I1(\rx_d[6] ), .O(\data_to_fifo[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3136.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3137 (.I0(rx_en_fifo), .I1(\rx_d[2] ), .O(\data_to_fifo[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3137.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3138 (.I0(rx_en_fifo), .I1(\rx_d[1] ), .O(\data_to_fifo[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3138.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3139 (.I0(n1751), .I1(n1749), .O(\i11/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3139.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3140 (.I0(\tx_dac_fsm_inst/sym_ctr[2] ), .I1(\tx_dac_fsm_inst/sym_ctr[3] ), 
            .O(n1633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3140.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3141 (.I0(n1633), .I1(\tx_dac_fsm_inst/sym_ctr[4] ), .O(n1753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3141.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3142 (.I0(n1753), .I1(\tx_dac_fsm_inst/sym_ctr[0] ), .O(\tx_dac_fsm_inst/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__3142.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__3143 (.I0(\tx_dac_fsm_inst/zctr[0] ), .I1(\tx_dac_fsm_inst/zctr[1] ), 
            .I2(\tx_dac_fsm_inst/zctr[2] ), .O(n1628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3143.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3144 (.I0(\tx_dac_fsm_inst/zctr[4] ), .I1(\tx_dac_fsm_inst/zctr[5] ), 
            .O(n1754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3144.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3145 (.I0(n1628), .I1(n1754), .I2(\tx_dac_fsm_inst/zctr[3] ), 
            .O(n1755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3145.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3146 (.I0(\tx_dac_fsm_inst/n283 ), .I1(\tx_dac_fsm_inst/n282 ), 
            .O(n1756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3146.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3147 (.I0(\tx_dac_fsm_inst/dctr[1]~FF_frt_1_q ), .I1(\tx_dac_fsm_inst/dctr[0] ), 
            .O(n1617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3147.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3148 (.I0(\tx_dac_fsm_inst/n280 ), .I1(\tx_dac_fsm_inst/n279 ), 
            .O(n1757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3148.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3149 (.I0(n1617), .I1(\tx_dac_fsm_inst/dctr[4]~FF_frt_0_q ), 
            .I2(\tx_dac_fsm_inst/dctr[3] ), .O(n1758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3149.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3150 (.I0(n1758), .I1(n1755), .I2(\tx_dac_fsm_inst/dac_config_reg[0] ), 
            .O(\tx_dac_fsm_inst/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__3150.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__3151 (.I0(\tx_dac_fsm_inst/n42 ), .I1(n1753), .O(\tx_dac_fsm_inst/n344 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3151.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3152 (.I0(\tx_dac_fsm_inst/dctr[1]~FF_frt_1_q ), .I1(\tx_dac_fsm_inst/dctr[3] ), 
            .I2(\tx_dac_fsm_inst/dctr[4]~FF_frt_0_q ), .O(n1759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3152.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3153 (.I0(\tx_dac_fsm_inst/dctr[0] ), .I1(\tx_dac_fsm_inst/dctr[2] ), 
            .I2(\tx_dac_fsm_inst/state_reg[2] ), .I3(n1759), .O(n1760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__3153.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__3154 (.I0(n1760), .I1(\tx_dac_fsm_inst/state_reg[0] ), 
            .I2(\tx_dac_fsm_inst/state_reg[2] ), .I3(n1754), .O(n1761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__3154.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__3155 (.I0(\tx_dac_fsm_inst/dac_config_reg[0] ), .I1(\tx_dac_fsm_inst/state_reg[2] ), 
            .I2(n1761), .O(n1762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__3155.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__3156 (.I0(\tx_dac_fsm_inst/dctr[3] ), .I1(\tx_dac_fsm_inst/dctr[1]~FF_frt_1_q ), 
            .I2(\tx_dac_fsm_inst/dctr[4]~FF_frt_0_q ), .I3(\tx_dac_fsm_inst/state_reg[0] ), 
            .O(n1763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__3156.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__3157 (.I0(n1763), .I1(\tx_dac_fsm_inst/state_reg[0] ), 
            .I2(\tx_dac_fsm_inst/state_reg[2] ), .I3(\tx_dac_fsm_inst/state_reg[3] ), 
            .O(n1764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfa3f */ ;
    defparam LUT__3157.LUTMASK = 16'hfa3f;
    EFX_LUT4 LUT__3158 (.I0(n1764), .I1(\tx_dac_fsm_inst/state_reg[1] ), 
            .O(n1438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3158.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3159 (.I0(\tx_dac_fsm_inst/sym_pos[2] ), .I1(\tx_dac_fsm_inst/sym_pos[1] ), 
            .I2(\tx_dac_fsm_inst/sym_pos[3] ), .I3(\tx_dac_fsm_inst/sym_pos[0] ), 
            .O(n1765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcf15 */ ;
    defparam LUT__3159.LUTMASK = 16'hcf15;
    EFX_LUT4 LUT__3160 (.I0(n1765), .I1(\tx_dac_fsm_inst/dac_config_reg[0] ), 
            .I2(\tx_dac_fsm_inst/state_reg[0] ), .I3(\tx_dac_fsm_inst/state_reg[1] ), 
            .O(n1766)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__3160.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__3161 (.I0(n1766), .I1(\tx_dac_fsm_inst/state_reg[2] ), 
            .I2(\tx_dac_fsm_inst/state_reg[3] ), .O(n1767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__3161.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__3162 (.I0(\tx_dac_fsm_inst/state_reg[1] ), .I1(n1762), 
            .I2(n1438), .I3(n1767), .O(n1410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3162.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3163 (.I0(\tx_dac_fsm_inst/state_reg[3] ), .I1(\tx_dac_fsm_inst/state_reg[0] ), 
            .I2(\tx_dac_fsm_inst/state_reg[1] ), .I3(\tx_dac_fsm_inst/state_reg[2] ), 
            .O(n1768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4110 */ ;
    defparam LUT__3163.LUTMASK = 16'h4110;
    EFX_LUT4 LUT__3164 (.I0(n1759), .I1(\tx_dac_fsm_inst/dac_config_reg[0] ), 
            .I2(\tx_dac_fsm_inst/state_reg[2] ), .I3(n1768), .O(n1411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacff */ ;
    defparam LUT__3164.LUTMASK = 16'hacff;
    EFX_LUT4 LUT__3165 (.I0(\tx_dac_fsm_inst/sym_ctr[1] ), .I1(n1159), .I2(n1753), 
            .O(\tx_dac_fsm_inst/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3165.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3166 (.I0(\tx_dac_fsm_inst/sym_ctr[2] ), .I1(n1156), .I2(n1753), 
            .O(\tx_dac_fsm_inst/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__3166.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__3167 (.I0(n1141), .I1(n1153), .I2(n1753), .O(\tx_dac_fsm_inst/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3167.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3168 (.I0(\tx_dac_fsm_inst/state_reg[0] ), .I1(\tx_dac_fsm_inst/state_reg[1] ), 
            .I2(\tx_dac_fsm_inst/state_reg[2] ), .I3(\tx_dac_fsm_inst/state_reg[3] ), 
            .O(n1415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__3168.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__3169 (.I0(\tx_dac_fsm_inst/state_reg[1] ), .I1(\tx_dac_fsm_inst/state_reg[2] ), 
            .O(n1769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3169.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3170 (.I0(n1769), .I1(\tx_dac_fsm_inst/state_reg[3] ), 
            .O(n1416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3170.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3171 (.I0(\tx_dac_fsm_inst/state_reg[3] ), .I1(\tx_dac_fsm_inst/state_reg[0] ), 
            .I2(n1769), .O(n1417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3171.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3172 (.I0(\tx_dac_fsm_inst/state_reg[2] ), .I1(\tx_dac_fsm_inst/state_reg[1] ), 
            .I2(\tx_dac_fsm_inst/state_reg[0] ), .O(n1418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3172.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3173 (.I0(\tx_dac_fsm_inst/zctr[0] ), .I1(n131), .O(\tx_dac_fsm_inst/n258 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3173.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3174 (.I0(n1139), .I1(n1150), .I2(n1753), .O(\tx_dac_fsm_inst/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3174.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3175 (.I0(\tx_dac_fsm_inst/dctr[0] ), .I1(n130), .O(\tx_dac_fsm_inst/n284 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3175.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3176 (.I0(n1710), .I1(n1744), .I2(\reg_addr[0] ), .O(rx_en_dac)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3176.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3177 (.I0(rx_en_dac), .I1(\rx_d[0] ), .O(data_to_dac)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3177.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3178 (.I0(\tx_dac_fsm_inst/sym_pos[0] ), .I1(\tx_dac_fsm_inst/sym_pos[1] ), 
            .O(\~tx_dac_fsm_inst/n431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3178.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3179 (.I0(\tx_dac_fsm_inst/sym_pos[0] ), .I1(\tx_dac_fsm_inst/sym_pos[1] ), 
            .I2(\tx_dac_fsm_inst/sym_pos[2] ), .O(\~tx_dac_fsm_inst/n436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3179.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3180 (.I0(\tx_dac_fsm_inst/sym_pos[0] ), .I1(\tx_dac_fsm_inst/sym_pos[1] ), 
            .I2(\tx_dac_fsm_inst/sym_pos[2] ), .I3(\tx_dac_fsm_inst/sym_pos[3] ), 
            .O(\~tx_dac_fsm_inst/n441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__3180.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__3181 (.I0(\tx_dac_fsm_inst/zctr[3] ), .I1(\tx_dac_fsm_inst/zctr[5] ), 
            .I2(\tx_dac_fsm_inst/zctr[4] ), .I3(\tx_dac_fsm_inst/state_reg[0] ), 
            .O(n1770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__3181.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__3182 (.I0(\tx_dac_fsm_inst/zctr[0] ), .I1(\tx_dac_fsm_inst/zctr[1] ), 
            .I2(\tx_dac_fsm_inst/zctr[2] ), .I3(\tx_dac_fsm_inst/dac_config_reg[0] ), 
            .O(n1771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3182.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3183 (.I0(n1769), .I1(n1770), .I2(n1771), .O(n1772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3183.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3184 (.I0(n1760), .I1(\tx_dac_fsm_inst/state_reg[0] ), 
            .I2(\tx_dac_fsm_inst/state_reg[1] ), .I3(n1772), .O(n1773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__3184.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__3185 (.I0(n1769), .I1(n1763), .I2(n1773), .I3(\tx_dac_fsm_inst/state_reg[3] ), 
            .O(n1436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h880f */ ;
    defparam LUT__3185.LUTMASK = 16'h880f;
    EFX_LUT4 LUT__3186 (.I0(\tx_dac_fsm_inst/state_reg[0] ), .I1(\tx_dac_fsm_inst/state_reg[2] ), 
            .I2(n1766), .I3(\tx_dac_fsm_inst/state_reg[3] ), .O(n1437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__3186.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__3187 (.I0(n1769), .I1(\tx_dac_fsm_inst/state_reg[3] ), 
            .I2(\tx_dac_fsm_inst/state_reg[0] ), .O(n1439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1818 */ ;
    defparam LUT__3187.LUTMASK = 16'h1818;
    EFX_LUT4 LUT__3188 (.I0(n131), .I1(n135), .O(\tx_dac_fsm_inst/n257 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3188.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3189 (.I0(n131), .I1(n1133), .O(\tx_dac_fsm_inst/n256 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3189.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3190 (.I0(n131), .I1(n1130), .O(\tx_dac_fsm_inst/n255 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3190.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3191 (.I0(n131), .I1(n1126), .O(\tx_dac_fsm_inst/n254 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3191.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3192 (.I0(n131), .I1(n1124), .O(\tx_dac_fsm_inst/n253 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3192.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3193 (.I0(n130), .I1(n138), .O(\tx_dac_fsm_inst/n283 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3193.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3194 (.I0(n130), .I1(n1118), .O(\tx_dac_fsm_inst/n282 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3194.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3195 (.I0(n130), .I1(n1095), .O(\tx_dac_fsm_inst/n281 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3195.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3196 (.I0(n130), .I1(n1092), .O(\tx_dac_fsm_inst/n280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3196.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3197 (.I0(n130), .I1(n1090), .O(\tx_dac_fsm_inst/n279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3197.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3198 (.I0(n1708), .I1(n1744), .I2(\reg_addr[0] ), .O(rx_en_fifo_length)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3198.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3199 (.I0(rx_en_fifo_length), .I1(\fifo_inst/wr_index[0] ), 
            .O(\fifo_inst/n153 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3199.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3200 (.I0(n1708), .I1(\reg_addr[0] ), .I2(n1744), .I3(n1745), 
            .O(ceg_net146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__3200.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__3201 (.I0(rx_en_fifo_length), .I1(\fifo_inst/rd_index[0] ), 
            .O(\fifo_inst/n162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3201.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3202 (.I0(\fifo_inst/wr_index[2] ), .I1(\fifo_inst/rd_index[2] ), 
            .I2(\fifo_inst/wr_index[3] ), .I3(\fifo_inst/rd_index[3] ), 
            .O(n1774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3202.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3203 (.I0(\fifo_inst/wr_index[0] ), .I1(\fifo_inst/rd_index[0] ), 
            .I2(\fifo_inst/wr_index[1] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3203.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3204 (.I0(\fifo_inst/wr_index[4] ), .I1(\fifo_inst/rd_index[4] ), 
            .I2(\fifo_inst/wr_index[5] ), .I3(\fifo_inst/rd_index[5] ), 
            .O(n1776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3204.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3205 (.I0(\fifo_inst/wr_index[6] ), .I1(\fifo_inst/rd_index[6] ), 
            .I2(\fifo_inst/wr_index[7] ), .I3(\fifo_inst/rd_index[7] ), 
            .O(n1777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3205.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3206 (.I0(n1774), .I1(n1775), .I2(n1776), .I3(n1777), 
            .O(n1778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3206.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3207 (.I0(\fifo_inst/sync_rd[0] ), .I1(n1745), .I2(\fifo_inst/sync_rd[1] ), 
            .I3(rx_en_fifo_length), .O(n1779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__3207.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__3208 (.I0(rx_en_fifo_length), .I1(n1778), .I2(n1779), 
            .O(ceg_net164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3208.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3209 (.I0(rx_en_fifo_length), .I1(\rx_d[0] ), .O(\data_to_fifo_length[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3209.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3210 (.I0(rx_en_fifo), .I1(n1745), .O(n1780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3210.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3211 (.I0(\i11/fifo_inst/buff[44][0] ), .I1(\i11/fifo_inst/buff[46][0] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__3211.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__3212 (.I0(\i11/fifo_inst/buff[47][0] ), .I1(\i11/fifo_inst/buff[45][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n1782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__3212.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__3213 (.I0(\i11/fifo_inst/buff[40][0] ), .I1(\i11/fifo_inst/buff[42][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3213.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3214 (.I0(\i11/fifo_inst/buff[43][0] ), .I1(\i11/fifo_inst/buff[41][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3214.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3215 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[1] ), 
            .I2(\fifo_inst/rd_index[2] ), .O(n1785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8787 */ ;
    defparam LUT__3215.LUTMASK = 16'h8787;
    EFX_LUT4 LUT__3216 (.I0(n1784), .I1(n1783), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1785), .O(n1786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3216.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3217 (.I0(n1782), .I1(n1781), .I2(n1786), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__3217.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__3218 (.I0(\i11/fifo_inst/buff[35][0] ), .I1(\i11/fifo_inst/buff[33][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3218.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3219 (.I0(\i11/fifo_inst/buff[32][0] ), .I1(\i11/fifo_inst/buff[34][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3219.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3220 (.I0(\i11/fifo_inst/buff[36][0] ), .I1(\i11/fifo_inst/buff[38][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3220.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3221 (.I0(\i11/fifo_inst/buff[39][0] ), .I1(\i11/fifo_inst/buff[37][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1790), .O(n1791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3221.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3222 (.I0(n1789), .I1(n1788), .I2(n1791), .I3(n1785), 
            .O(n1792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3222.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3223 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[1] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[3] ), 
            .O(n1793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3223.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3224 (.I0(n1793), .I1(\fifo_inst/rd_index[4] ), .I2(\fifo_inst/rd_index[5] ), 
            .O(n1794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7e7 */ ;
    defparam LUT__3224.LUTMASK = 16'he7e7;
    EFX_LUT4 LUT__3225 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[1] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[3] ), 
            .O(n1795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h807f */ ;
    defparam LUT__3225.LUTMASK = 16'h807f;
    EFX_LUT4 LUT__3226 (.I0(n1792), .I1(n1787), .I2(n1794), .I3(n1795), 
            .O(n1796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3226.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3227 (.I0(\i11/fifo_inst/buff[28][0] ), .I1(\i11/fifo_inst/buff[30][0] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__3227.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__3228 (.I0(\i11/fifo_inst/buff[31][0] ), .I1(\i11/fifo_inst/buff[29][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n1798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__3228.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__3229 (.I0(\i11/fifo_inst/buff[24][0] ), .I1(\i11/fifo_inst/buff[26][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3229.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3230 (.I0(\i11/fifo_inst/buff[27][0] ), .I1(\i11/fifo_inst/buff[25][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3230.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3231 (.I0(n1800), .I1(n1799), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1785), .O(n1801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3231.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3232 (.I0(n1798), .I1(n1797), .I2(n1801), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__3232.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__3233 (.I0(\i11/fifo_inst/buff[19][0] ), .I1(\i11/fifo_inst/buff[17][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3233.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3234 (.I0(\i11/fifo_inst/buff[16][0] ), .I1(\i11/fifo_inst/buff[18][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3234.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3235 (.I0(\i11/fifo_inst/buff[20][0] ), .I1(\i11/fifo_inst/buff[22][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3235.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3236 (.I0(\i11/fifo_inst/buff[23][0] ), .I1(\i11/fifo_inst/buff[21][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1805), .O(n1806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3236.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3237 (.I0(n1804), .I1(n1803), .I2(n1806), .I3(n1785), 
            .O(n1807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3237.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3238 (.I0(\fifo_inst/rd_index[5] ), .I1(n1793), .I2(\fifo_inst/rd_index[4] ), 
            .O(n1808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3238.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__3239 (.I0(n1807), .I1(n1802), .I2(n1795), .I3(n1808), 
            .O(n1809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3239.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3240 (.I0(\i11/fifo_inst/buff[52][0] ), .I1(\i11/fifo_inst/buff[54][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3240.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3241 (.I0(\i11/fifo_inst/buff[53][0] ), .I1(\i11/fifo_inst/buff[55][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1810), .O(n1811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__3241.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__3242 (.I0(\i11/fifo_inst/buff[48][0] ), .I1(\i11/fifo_inst/buff[50][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3242.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3243 (.I0(\i11/fifo_inst/buff[51][0] ), .I1(\i11/fifo_inst/buff[49][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1812), .O(n1813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3243.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3244 (.I0(n1813), .I1(n1811), .I2(n1785), .I3(n1795), 
            .O(n1814)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha300 */ ;
    defparam LUT__3244.LUTMASK = 16'ha300;
    EFX_LUT4 LUT__3245 (.I0(\i11/fifo_inst/buff[2][0] ), .I1(\i11/fifo_inst/buff[0][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3245.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3246 (.I0(\i11/fifo_inst/buff[3][0] ), .I1(\i11/fifo_inst/buff[1][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3246.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3247 (.I0(n1816), .I1(n1815), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1785), .O(n1817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3247.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3248 (.I0(\i11/fifo_inst/buff[6][0] ), .I1(\i11/fifo_inst/buff[4][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n1818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__3248.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__3249 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[2] ), 
            .O(n1819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3249.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3250 (.I0(\i11/fifo_inst/buff[7][0] ), .I1(\i11/fifo_inst/buff[5][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3250.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3251 (.I0(n1820), .I1(n1819), .I2(n1818), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__3251.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__3252 (.I0(n1793), .I1(\fifo_inst/rd_index[4] ), .I2(\fifo_inst/rd_index[5] ), 
            .O(n1822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7e7e */ ;
    defparam LUT__3252.LUTMASK = 16'h7e7e;
    EFX_LUT4 LUT__3253 (.I0(n1817), .I1(n1821), .I2(n1795), .I3(n1822), 
            .O(n1823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__3253.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__3254 (.I0(\i11/fifo_inst/buff[63][0] ), .I1(\i11/fifo_inst/buff[61][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n1824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__3254.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__3255 (.I0(\i11/fifo_inst/buff[60][0] ), .I1(\i11/fifo_inst/buff[62][0] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__3255.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__3256 (.I0(n1824), .I1(n1825), .I2(n1795), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__3256.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__3257 (.I0(\i11/fifo_inst/buff[56][0] ), .I1(\i11/fifo_inst/buff[58][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3257.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3258 (.I0(\i11/fifo_inst/buff[59][0] ), .I1(\i11/fifo_inst/buff[57][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1827), .O(n1828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3258.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3259 (.I0(n1793), .I1(\fifo_inst/rd_index[4] ), .I2(\fifo_inst/rd_index[5] ), 
            .O(n1829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__3259.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__3260 (.I0(n1828), .I1(n1785), .I2(n1826), .I3(n1829), 
            .O(n1830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__3260.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__3261 (.I0(\i11/fifo_inst/buff[12][0] ), .I1(\i11/fifo_inst/buff[14][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3261.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3262 (.I0(\i11/fifo_inst/buff[13][0] ), .I1(\i11/fifo_inst/buff[15][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1831), .O(n1832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__3262.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__3263 (.I0(\i11/fifo_inst/buff[8][0] ), .I1(\i11/fifo_inst/buff[10][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3263.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3264 (.I0(\i11/fifo_inst/buff[11][0] ), .I1(\i11/fifo_inst/buff[9][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1833), .O(n1834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3264.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3265 (.I0(n1834), .I1(n1832), .I2(n1795), .I3(n1785), 
            .O(n1835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__3265.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__3266 (.I0(n1835), .I1(n1823), .I2(n1814), .I3(n1830), 
            .O(n1836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__3266.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__3267 (.I0(n1793), .I1(\fifo_inst/rd_index[4] ), .I2(\fifo_inst/rd_index[5] ), 
            .I3(\fifo_inst/rd_index[6] ), .O(n1837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h807f */ ;
    defparam LUT__3267.LUTMASK = 16'h807f;
    EFX_LUT4 LUT__3268 (.I0(n1778), .I1(n1837), .I2(ceg_net146), .O(n1838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3268.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3269 (.I0(n1809), .I1(n1796), .I2(n1836), .I3(n1838), 
            .O(n1839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__3269.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__3270 (.I0(\i11/fifo_inst/buff[115][0] ), .I1(\i11/fifo_inst/buff[113][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3270.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3271 (.I0(\i11/fifo_inst/buff[112][0] ), .I1(\i11/fifo_inst/buff[114][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3271.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3272 (.I0(\i11/fifo_inst/buff[116][0] ), .I1(\i11/fifo_inst/buff[118][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3272.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3273 (.I0(\i11/fifo_inst/buff[119][0] ), .I1(\i11/fifo_inst/buff[117][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1842), .O(n1843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3273.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3274 (.I0(n1841), .I1(n1840), .I2(n1843), .I3(n1785), 
            .O(n1844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3274.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3275 (.I0(\i11/fifo_inst/buff[123][0] ), .I1(\i11/fifo_inst/buff[121][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3275.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3276 (.I0(\i11/fifo_inst/buff[120][0] ), .I1(\i11/fifo_inst/buff[122][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3276.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3277 (.I0(\i11/fifo_inst/buff[124][0] ), .I1(\i11/fifo_inst/buff[126][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3277.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3278 (.I0(\i11/fifo_inst/buff[127][0] ), .I1(\i11/fifo_inst/buff[125][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1847), .O(n1848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3278.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3279 (.I0(n1846), .I1(n1845), .I2(n1848), .I3(n1785), 
            .O(n1849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3279.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3280 (.I0(n1849), .I1(n1844), .I2(n1795), .I3(n1829), 
            .O(n1850)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3280.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3281 (.I0(\i11/fifo_inst/buff[76][0] ), .I1(\i11/fifo_inst/buff[78][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3281.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3282 (.I0(\i11/fifo_inst/buff[79][0] ), .I1(\i11/fifo_inst/buff[77][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3282.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3283 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[1] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[3] ), 
            .O(n1853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__3283.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__3284 (.I0(n1852), .I1(n1851), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1853), .O(n1854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3284.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3285 (.I0(\i11/fifo_inst/buff[64][0] ), .I1(\i11/fifo_inst/buff[66][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3285.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3286 (.I0(\i11/fifo_inst/buff[67][0] ), .I1(\i11/fifo_inst/buff[65][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3286.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3287 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[1] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[3] ), 
            .O(n1857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ff8 */ ;
    defparam LUT__3287.LUTMASK = 16'h7ff8;
    EFX_LUT4 LUT__3288 (.I0(n1856), .I1(n1855), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3288.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3289 (.I0(\i11/fifo_inst/buff[68][0] ), .I1(\i11/fifo_inst/buff[70][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3289.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3290 (.I0(\i11/fifo_inst/buff[71][0] ), .I1(\i11/fifo_inst/buff[69][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3290.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3291 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[1] ), 
            .I2(\fifo_inst/rd_index[3] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n1861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__3291.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__3292 (.I0(n1860), .I1(n1859), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n1862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3292.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3293 (.I0(\i11/fifo_inst/buff[72][0] ), .I1(\i11/fifo_inst/buff[74][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3293.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3294 (.I0(\i11/fifo_inst/buff[75][0] ), .I1(\i11/fifo_inst/buff[73][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3294.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3295 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[1] ), 
            .I2(\fifo_inst/rd_index[3] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n1865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf78f */ ;
    defparam LUT__3295.LUTMASK = 16'hf78f;
    EFX_LUT4 LUT__3296 (.I0(n1864), .I1(n1863), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3296.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3297 (.I0(n1854), .I1(n1858), .I2(n1862), .I3(n1866), 
            .O(n1867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3297.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3298 (.I0(\i11/fifo_inst/buff[80][0] ), .I1(\i11/fifo_inst/buff[82][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3298.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3299 (.I0(\i11/fifo_inst/buff[83][0] ), .I1(\i11/fifo_inst/buff[81][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3299.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3300 (.I0(n1869), .I1(n1868), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3300.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3301 (.I0(\i11/fifo_inst/buff[92][0] ), .I1(\i11/fifo_inst/buff[94][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3301.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3302 (.I0(\i11/fifo_inst/buff[95][0] ), .I1(\i11/fifo_inst/buff[93][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3302.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3303 (.I0(n1872), .I1(n1871), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1853), .O(n1873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3303.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3304 (.I0(\i11/fifo_inst/buff[88][0] ), .I1(\i11/fifo_inst/buff[90][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3304.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3305 (.I0(\i11/fifo_inst/buff[91][0] ), .I1(\i11/fifo_inst/buff[89][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3305.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3306 (.I0(n1875), .I1(n1874), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3306.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3307 (.I0(\i11/fifo_inst/buff[84][0] ), .I1(\i11/fifo_inst/buff[86][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3307.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3308 (.I0(\i11/fifo_inst/buff[87][0] ), .I1(\i11/fifo_inst/buff[85][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3308.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3309 (.I0(n1878), .I1(n1877), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n1879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3309.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3310 (.I0(n1870), .I1(n1873), .I2(n1876), .I3(n1879), 
            .O(n1880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3310.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3311 (.I0(n1793), .I1(\fifo_inst/rd_index[4] ), .I2(\fifo_inst/rd_index[5] ), 
            .O(n1881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8787 */ ;
    defparam LUT__3311.LUTMASK = 16'h8787;
    EFX_LUT4 LUT__3312 (.I0(n1793), .I1(\fifo_inst/rd_index[4] ), .O(n1882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__3312.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__3313 (.I0(n1880), .I1(n1867), .I2(n1882), .I3(n1881), 
            .O(n1883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3313.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3314 (.I0(\i11/fifo_inst/buff[99][0] ), .I1(\i11/fifo_inst/buff[97][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3314.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3315 (.I0(\i11/fifo_inst/buff[96][0] ), .I1(\i11/fifo_inst/buff[98][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3315.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3316 (.I0(\i11/fifo_inst/buff[100][0] ), .I1(\i11/fifo_inst/buff[102][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3316.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3317 (.I0(\i11/fifo_inst/buff[103][0] ), .I1(\i11/fifo_inst/buff[101][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1886), .O(n1887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3317.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3318 (.I0(n1885), .I1(n1884), .I2(n1887), .I3(n1785), 
            .O(n1888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3318.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3319 (.I0(\i11/fifo_inst/buff[107][0] ), .I1(\i11/fifo_inst/buff[105][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3319.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3320 (.I0(\i11/fifo_inst/buff[104][0] ), .I1(\i11/fifo_inst/buff[106][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3320.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3321 (.I0(\i11/fifo_inst/buff[108][0] ), .I1(\i11/fifo_inst/buff[110][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3321.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3322 (.I0(\i11/fifo_inst/buff[111][0] ), .I1(\i11/fifo_inst/buff[109][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1891), .O(n1892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3322.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3323 (.I0(n1890), .I1(n1889), .I2(n1892), .I3(n1785), 
            .O(n1893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3323.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3324 (.I0(n1893), .I1(n1888), .I2(n1794), .I3(n1795), 
            .O(n1894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3324.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3325 (.I0(n1778), .I1(n1837), .I2(ceg_net146), .O(n1895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3325.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3326 (.I0(n1883), .I1(n1894), .I2(n1850), .I3(n1895), 
            .O(n1896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__3326.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__3327 (.I0(n1780), .I1(\rx_d[0] ), .I2(n1839), .I3(n1896), 
            .O(\fifo_inst/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__3327.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__3328 (.I0(n1778), .I1(n1745), .I2(n1779), .O(ceg_net242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3328.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3329 (.I0(rx_en_fifo_length), .I1(n141), .O(\fifo_inst/n152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3329.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3330 (.I0(rx_en_fifo_length), .I1(n1083), .O(\fifo_inst/n151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3330.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3331 (.I0(rx_en_fifo_length), .I1(n1080), .O(\fifo_inst/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3331.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3332 (.I0(rx_en_fifo_length), .I1(n1077), .O(\fifo_inst/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3332.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3333 (.I0(rx_en_fifo_length), .I1(n1073), .O(\fifo_inst/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3333.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3334 (.I0(rx_en_fifo_length), .I1(n1070), .O(\fifo_inst/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3334.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3335 (.I0(rx_en_fifo_length), .I1(n1067), .O(\fifo_inst/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3335.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3336 (.I0(rx_en_fifo_length), .I1(\fifo_inst/rd_index[0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(\fifo_inst/n161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3336.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__3337 (.I0(rx_en_fifo_length), .I1(n1785), .O(\fifo_inst/n160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3337.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3338 (.I0(rx_en_fifo_length), .I1(n1795), .O(\fifo_inst/n159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3338.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3339 (.I0(rx_en_fifo_length), .I1(n1882), .O(\fifo_inst/n158 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3339.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3340 (.I0(rx_en_fifo_length), .I1(n1881), .O(\fifo_inst/n157 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3340.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3341 (.I0(rx_en_fifo_length), .I1(n1837), .O(\fifo_inst/n156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3341.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3342 (.I0(n1837), .I1(\fifo_inst/rd_index[6] ), .I2(rx_en_fifo_length), 
            .I3(\fifo_inst/rd_index[7] ), .O(\fifo_inst/n155 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__3342.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__3343 (.I0(rx_en_fifo_length), .I1(\rx_d[1] ), .O(\data_to_fifo_length[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3343.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3344 (.I0(rx_en_fifo_length), .I1(\rx_d[2] ), .O(\data_to_fifo_length[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3344.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3345 (.I0(rx_en_fifo_length), .I1(\rx_d[3] ), .O(\data_to_fifo_length[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3345.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3346 (.I0(rx_en_fifo_length), .I1(\rx_d[4] ), .O(\data_to_fifo_length[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3346.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3347 (.I0(rx_en_fifo_length), .I1(\rx_d[5] ), .O(\data_to_fifo_length[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3347.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3348 (.I0(rx_en_fifo_length), .I1(\rx_d[6] ), .O(\data_to_fifo_length[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3348.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3349 (.I0(rx_en_fifo_length), .I1(\rx_d[7] ), .O(\data_to_fifo_length[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3349.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3350 (.I0(n1747), .I1(n1752), .O(\i11/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3350.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3351 (.I0(\i11/fifo_inst/buff[87][1] ), .I1(\i11/fifo_inst/buff[85][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3351.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3352 (.I0(\i11/fifo_inst/buff[84][1] ), .I1(\i11/fifo_inst/buff[86][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3352.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3353 (.I0(\i11/fifo_inst/buff[116][1] ), .I1(\i11/fifo_inst/buff[118][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3353.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3354 (.I0(\i11/fifo_inst/buff[119][1] ), .I1(\i11/fifo_inst/buff[117][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1899), .O(n1900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3354.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3355 (.I0(n1898), .I1(n1897), .I2(n1900), .I3(n1881), 
            .O(n1901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3355.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3356 (.I0(\i11/fifo_inst/buff[83][1] ), .I1(\i11/fifo_inst/buff[81][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3356.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3357 (.I0(\i11/fifo_inst/buff[80][1] ), .I1(\i11/fifo_inst/buff[82][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3357.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3358 (.I0(\i11/fifo_inst/buff[112][1] ), .I1(\i11/fifo_inst/buff[114][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3358.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3359 (.I0(\i11/fifo_inst/buff[115][1] ), .I1(\i11/fifo_inst/buff[113][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1904), .O(n1905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3359.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3360 (.I0(n1903), .I1(n1902), .I2(n1905), .I3(n1881), 
            .O(n1906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3360.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3361 (.I0(n1906), .I1(n1901), .I2(n1785), .I3(n1795), 
            .O(n1907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__3361.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__3362 (.I0(\i11/fifo_inst/buff[95][1] ), .I1(\i11/fifo_inst/buff[93][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3362.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3363 (.I0(\i11/fifo_inst/buff[92][1] ), .I1(\i11/fifo_inst/buff[94][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3363.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3364 (.I0(\i11/fifo_inst/buff[91][1] ), .I1(\i11/fifo_inst/buff[89][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3364.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3365 (.I0(\i11/fifo_inst/buff[88][1] ), .I1(\i11/fifo_inst/buff[90][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3365.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3366 (.I0(n1911), .I1(n1910), .I2(n1785), .I3(\fifo_inst/rd_index[5] ), 
            .O(n1912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__3366.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__3367 (.I0(n1909), .I1(n1785), .I2(n1908), .I3(n1912), 
            .O(n1913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__3367.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__3368 (.I0(\i11/fifo_inst/buff[124][1] ), .I1(\i11/fifo_inst/buff[126][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3368.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3369 (.I0(\i11/fifo_inst/buff[127][1] ), .I1(\i11/fifo_inst/buff[125][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1914), .O(n1915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3369.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3370 (.I0(\i11/fifo_inst/buff[120][1] ), .I1(\i11/fifo_inst/buff[122][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3370.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3371 (.I0(\i11/fifo_inst/buff[123][1] ), .I1(\i11/fifo_inst/buff[121][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1916), .O(n1917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3371.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3372 (.I0(n1917), .I1(n1915), .I2(n1785), .I3(\fifo_inst/rd_index[5] ), 
            .O(n1918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3372.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3373 (.I0(n1918), .I1(n1913), .I2(n1795), .I3(n1882), 
            .O(n1919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f1 */ ;
    defparam LUT__3373.LUTMASK = 16'h00f1;
    EFX_LUT4 LUT__3374 (.I0(\i11/fifo_inst/buff[68][1] ), .I1(\i11/fifo_inst/buff[70][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3374.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3375 (.I0(\i11/fifo_inst/buff[71][1] ), .I1(\i11/fifo_inst/buff[69][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3375.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3376 (.I0(n1921), .I1(n1920), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n1922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3376.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3377 (.I0(\i11/fifo_inst/buff[76][1] ), .I1(\i11/fifo_inst/buff[78][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3377.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3378 (.I0(\i11/fifo_inst/buff[79][1] ), .I1(\i11/fifo_inst/buff[77][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3378.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3379 (.I0(n1924), .I1(n1923), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1853), .O(n1925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3379.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3380 (.I0(\i11/fifo_inst/buff[64][1] ), .I1(\i11/fifo_inst/buff[66][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3380.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3381 (.I0(\i11/fifo_inst/buff[67][1] ), .I1(\i11/fifo_inst/buff[65][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3381.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3382 (.I0(n1927), .I1(n1926), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3382.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3383 (.I0(\i11/fifo_inst/buff[72][1] ), .I1(\i11/fifo_inst/buff[74][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3383.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3384 (.I0(\i11/fifo_inst/buff[75][1] ), .I1(\i11/fifo_inst/buff[73][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3384.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3385 (.I0(n1930), .I1(n1929), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3385.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3386 (.I0(n1922), .I1(n1925), .I2(n1928), .I3(n1931), 
            .O(n1932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3386.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3387 (.I0(\i11/fifo_inst/buff[96][1] ), .I1(\i11/fifo_inst/buff[98][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3387.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3388 (.I0(\i11/fifo_inst/buff[99][1] ), .I1(\i11/fifo_inst/buff[97][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3388.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3389 (.I0(n1934), .I1(n1933), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3389.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3390 (.I0(\i11/fifo_inst/buff[108][1] ), .I1(\i11/fifo_inst/buff[110][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3390.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3391 (.I0(\i11/fifo_inst/buff[111][1] ), .I1(\i11/fifo_inst/buff[109][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3391.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3392 (.I0(n1937), .I1(n1936), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1853), .O(n1938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3392.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3393 (.I0(\i11/fifo_inst/buff[100][1] ), .I1(\i11/fifo_inst/buff[102][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3393.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3394 (.I0(\i11/fifo_inst/buff[103][1] ), .I1(\i11/fifo_inst/buff[101][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3394.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3395 (.I0(n1940), .I1(n1939), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n1941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3395.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3396 (.I0(\i11/fifo_inst/buff[104][1] ), .I1(\i11/fifo_inst/buff[106][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3396.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3397 (.I0(\i11/fifo_inst/buff[107][1] ), .I1(\i11/fifo_inst/buff[105][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n1943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3397.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3398 (.I0(n1943), .I1(n1942), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3398.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3399 (.I0(n1935), .I1(n1938), .I2(n1941), .I3(n1944), 
            .O(n1945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3399.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3400 (.I0(n1945), .I1(n1932), .I2(n1881), .I3(n1882), 
            .O(n1946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3400.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3401 (.I0(n1907), .I1(n1919), .I2(n1946), .I3(n1895), 
            .O(n1947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__3401.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__3402 (.I0(\i11/fifo_inst/buff[14][1] ), .I1(\i11/fifo_inst/buff[12][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n1948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__3402.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__3403 (.I0(n1948), .I1(\fifo_inst/rd_index[0] ), .O(n1949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3403.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3404 (.I0(\i11/fifo_inst/buff[8][1] ), .I1(\i11/fifo_inst/buff[10][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3404.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3405 (.I0(\i11/fifo_inst/buff[11][1] ), .I1(\i11/fifo_inst/buff[9][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1950), .O(n1951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3405.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3406 (.I0(\i11/fifo_inst/buff[13][1] ), .I1(\i11/fifo_inst/buff[15][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(n1819), .O(n1952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__3406.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__3407 (.I0(n1785), .I1(n1951), .I2(n1952), .I3(n1949), 
            .O(n1953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__3407.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__3408 (.I0(\i11/fifo_inst/buff[3][1] ), .I1(\i11/fifo_inst/buff[1][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3408.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3409 (.I0(\i11/fifo_inst/buff[2][1] ), .I1(\i11/fifo_inst/buff[0][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3409.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3410 (.I0(\i11/fifo_inst/buff[4][1] ), .I1(\i11/fifo_inst/buff[6][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3410.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3411 (.I0(\i11/fifo_inst/buff[7][1] ), .I1(\i11/fifo_inst/buff[5][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1956), .O(n1957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3411.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3412 (.I0(n1955), .I1(n1954), .I2(n1957), .I3(n1785), 
            .O(n1958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3412.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3413 (.I0(n1958), .I1(n1953), .I2(n1822), .I3(n1795), 
            .O(n1959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3413.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3414 (.I0(\i11/fifo_inst/buff[22][1] ), .I1(\i11/fifo_inst/buff[20][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n1960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__3414.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__3415 (.I0(n1960), .I1(\fifo_inst/rd_index[0] ), .O(n1961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3415.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3416 (.I0(\i11/fifo_inst/buff[16][1] ), .I1(\i11/fifo_inst/buff[18][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3416.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3417 (.I0(\i11/fifo_inst/buff[19][1] ), .I1(\i11/fifo_inst/buff[17][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1962), .O(n1963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3417.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3418 (.I0(\i11/fifo_inst/buff[21][1] ), .I1(\i11/fifo_inst/buff[23][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(n1819), .O(n1964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__3418.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__3419 (.I0(n1785), .I1(n1963), .I2(n1964), .I3(n1961), 
            .O(n1965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__3419.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__3420 (.I0(\i11/fifo_inst/buff[27][1] ), .I1(\i11/fifo_inst/buff[25][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3420.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3421 (.I0(\i11/fifo_inst/buff[24][1] ), .I1(\i11/fifo_inst/buff[26][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3421.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3422 (.I0(\i11/fifo_inst/buff[28][1] ), .I1(\i11/fifo_inst/buff[30][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3422.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3423 (.I0(\i11/fifo_inst/buff[31][1] ), .I1(\i11/fifo_inst/buff[29][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1968), .O(n1969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3423.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3424 (.I0(n1967), .I1(n1966), .I2(n1969), .I3(n1785), 
            .O(n1970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3424.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3425 (.I0(n1970), .I1(n1965), .I2(n1795), .I3(n1808), 
            .O(n1971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3425.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3426 (.I0(\i11/fifo_inst/buff[44][1] ), .I1(\i11/fifo_inst/buff[46][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3426.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3427 (.I0(\i11/fifo_inst/buff[45][1] ), .I1(\i11/fifo_inst/buff[47][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1972), .O(n1973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__3427.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__3428 (.I0(\i11/fifo_inst/buff[40][1] ), .I1(\i11/fifo_inst/buff[42][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3428.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3429 (.I0(\i11/fifo_inst/buff[43][1] ), .I1(\i11/fifo_inst/buff[41][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1974), .O(n1975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3429.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3430 (.I0(n1975), .I1(n1973), .I2(n1795), .I3(n1785), 
            .O(n1976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__3430.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__3431 (.I0(\i11/fifo_inst/buff[39][1] ), .I1(\i11/fifo_inst/buff[37][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n1977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__3431.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__3432 (.I0(\i11/fifo_inst/buff[36][1] ), .I1(\i11/fifo_inst/buff[38][1] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__3432.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__3433 (.I0(n1977), .I1(n1978), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1795), .O(n1979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;
    defparam LUT__3433.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__3434 (.I0(\i11/fifo_inst/buff[32][1] ), .I1(\i11/fifo_inst/buff[34][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3434.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3435 (.I0(\i11/fifo_inst/buff[35][1] ), .I1(\i11/fifo_inst/buff[33][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1980), .O(n1981)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3435.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3436 (.I0(n1981), .I1(n1785), .I2(n1979), .I3(n1794), 
            .O(n1982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__3436.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__3437 (.I0(\i11/fifo_inst/buff[52][1] ), .I1(\i11/fifo_inst/buff[54][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3437.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3438 (.I0(\i11/fifo_inst/buff[53][1] ), .I1(\i11/fifo_inst/buff[55][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1983), .O(n1984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__3438.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__3439 (.I0(\i11/fifo_inst/buff[48][1] ), .I1(\i11/fifo_inst/buff[50][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3439.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3440 (.I0(\i11/fifo_inst/buff[51][1] ), .I1(\i11/fifo_inst/buff[49][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1985), .O(n1986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3440.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3441 (.I0(n1986), .I1(n1984), .I2(n1785), .I3(n1795), 
            .O(n1987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha300 */ ;
    defparam LUT__3441.LUTMASK = 16'ha300;
    EFX_LUT4 LUT__3442 (.I0(\i11/fifo_inst/buff[63][1] ), .I1(\i11/fifo_inst/buff[61][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n1988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__3442.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__3443 (.I0(\i11/fifo_inst/buff[60][1] ), .I1(\i11/fifo_inst/buff[62][1] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__3443.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__3444 (.I0(n1988), .I1(n1989), .I2(n1795), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__3444.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__3445 (.I0(\i11/fifo_inst/buff[56][1] ), .I1(\i11/fifo_inst/buff[58][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3445.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3446 (.I0(\i11/fifo_inst/buff[59][1] ), .I1(\i11/fifo_inst/buff[57][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1991), .O(n1992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3446.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3447 (.I0(n1992), .I1(n1785), .I2(n1990), .I3(n1829), 
            .O(n1993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__3447.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__3448 (.I0(n1987), .I1(n1993), .I2(n1976), .I3(n1982), 
            .O(n1994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__3448.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__3449 (.I0(n1971), .I1(n1959), .I2(n1994), .I3(n1838), 
            .O(n1995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__3449.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__3450 (.I0(n1780), .I1(\rx_d[1] ), .I2(n1947), .I3(n1995), 
            .O(\fifo_inst/n143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__3450.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__3451 (.I0(\i11/fifo_inst/buff[55][2] ), .I1(\i11/fifo_inst/buff[53][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3451.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3452 (.I0(\i11/fifo_inst/buff[52][2] ), .I1(\i11/fifo_inst/buff[54][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n1997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3452.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3453 (.I0(\i11/fifo_inst/buff[48][2] ), .I1(\i11/fifo_inst/buff[50][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n1998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3453.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3454 (.I0(\i11/fifo_inst/buff[51][2] ), .I1(\i11/fifo_inst/buff[49][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n1998), .O(n1999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3454.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3455 (.I0(n1997), .I1(n1996), .I2(n1999), .I3(n1785), 
            .O(n2000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__3455.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__3456 (.I0(\i11/fifo_inst/buff[59][2] ), .I1(\i11/fifo_inst/buff[57][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3456.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3457 (.I0(\i11/fifo_inst/buff[56][2] ), .I1(\i11/fifo_inst/buff[58][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3457.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3458 (.I0(\i11/fifo_inst/buff[60][2] ), .I1(\i11/fifo_inst/buff[62][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3458.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3459 (.I0(\i11/fifo_inst/buff[63][2] ), .I1(\i11/fifo_inst/buff[61][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2003), .O(n2004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3459.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3460 (.I0(n2002), .I1(n2001), .I2(n2004), .I3(n1785), 
            .O(n2005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3460.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3461 (.I0(n2005), .I1(n2000), .I2(n1795), .I3(n1829), 
            .O(n2006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3461.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3462 (.I0(\i11/fifo_inst/buff[35][2] ), .I1(\i11/fifo_inst/buff[33][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3462.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3463 (.I0(\i11/fifo_inst/buff[32][2] ), .I1(\i11/fifo_inst/buff[34][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3463.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3464 (.I0(\i11/fifo_inst/buff[36][2] ), .I1(\i11/fifo_inst/buff[38][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3464.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3465 (.I0(\i11/fifo_inst/buff[39][2] ), .I1(\i11/fifo_inst/buff[37][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2009), .O(n2010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3465.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3466 (.I0(n2008), .I1(n2007), .I2(n2010), .I3(n1785), 
            .O(n2011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3466.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3467 (.I0(\i11/fifo_inst/buff[43][2] ), .I1(\i11/fifo_inst/buff[41][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3467.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3468 (.I0(\i11/fifo_inst/buff[40][2] ), .I1(\i11/fifo_inst/buff[42][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3468.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3469 (.I0(\i11/fifo_inst/buff[44][2] ), .I1(\i11/fifo_inst/buff[46][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3469.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3470 (.I0(\i11/fifo_inst/buff[47][2] ), .I1(\i11/fifo_inst/buff[45][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2014), .O(n2015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3470.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3471 (.I0(n2013), .I1(n2012), .I2(n2015), .I3(n1785), 
            .O(n2016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3471.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3472 (.I0(n2016), .I1(n2011), .I2(n1794), .I3(n1795), 
            .O(n2017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3472.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3473 (.I0(\i11/fifo_inst/buff[3][2] ), .I1(\i11/fifo_inst/buff[1][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3473.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3474 (.I0(\i11/fifo_inst/buff[2][2] ), .I1(\i11/fifo_inst/buff[0][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3474.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3475 (.I0(\i11/fifo_inst/buff[4][2] ), .I1(\i11/fifo_inst/buff[6][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3475.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3476 (.I0(\i11/fifo_inst/buff[7][2] ), .I1(\i11/fifo_inst/buff[5][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2020), .O(n2021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3476.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3477 (.I0(n2019), .I1(n2018), .I2(n2021), .I3(n1785), 
            .O(n2022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3477.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3478 (.I0(\i11/fifo_inst/buff[11][2] ), .I1(\i11/fifo_inst/buff[9][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3478.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3479 (.I0(\i11/fifo_inst/buff[8][2] ), .I1(\i11/fifo_inst/buff[10][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3479.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3480 (.I0(\i11/fifo_inst/buff[12][2] ), .I1(\i11/fifo_inst/buff[14][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3480.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3481 (.I0(\i11/fifo_inst/buff[15][2] ), .I1(\i11/fifo_inst/buff[13][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2025), .O(n2026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3481.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3482 (.I0(n2024), .I1(n2023), .I2(n2026), .I3(n1785), 
            .O(n2027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3482.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3483 (.I0(n2027), .I1(n2022), .I2(n1822), .I3(n1795), 
            .O(n2028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3483.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3484 (.I0(\i11/fifo_inst/buff[19][2] ), .I1(\i11/fifo_inst/buff[17][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3484.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3485 (.I0(\i11/fifo_inst/buff[16][2] ), .I1(\i11/fifo_inst/buff[18][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3485.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3486 (.I0(\i11/fifo_inst/buff[20][2] ), .I1(\i11/fifo_inst/buff[22][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3486.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3487 (.I0(\i11/fifo_inst/buff[23][2] ), .I1(\i11/fifo_inst/buff[21][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2031), .O(n2032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3487.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3488 (.I0(n2030), .I1(n2029), .I2(n2032), .I3(n1785), 
            .O(n2033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3488.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3489 (.I0(\i11/fifo_inst/buff[27][2] ), .I1(\i11/fifo_inst/buff[25][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3489.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3490 (.I0(\i11/fifo_inst/buff[24][2] ), .I1(\i11/fifo_inst/buff[26][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3490.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3491 (.I0(\i11/fifo_inst/buff[28][2] ), .I1(\i11/fifo_inst/buff[30][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3491.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3492 (.I0(\i11/fifo_inst/buff[31][2] ), .I1(\i11/fifo_inst/buff[29][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2036), .O(n2037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3492.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3493 (.I0(n2035), .I1(n2034), .I2(n2037), .I3(n1785), 
            .O(n2038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3493.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3494 (.I0(n2038), .I1(n2033), .I2(n1795), .I3(n1808), 
            .O(n2039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3494.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3495 (.I0(n2006), .I1(n2017), .I2(n2028), .I3(n2039), 
            .O(n2040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3495.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3496 (.I0(\i11/fifo_inst/buff[116][2] ), .I1(\i11/fifo_inst/buff[118][2] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__3496.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__3497 (.I0(\i11/fifo_inst/buff[119][2] ), .I1(\i11/fifo_inst/buff[117][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n2042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__3497.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__3498 (.I0(\i11/fifo_inst/buff[112][2] ), .I1(\i11/fifo_inst/buff[114][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3498.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3499 (.I0(\i11/fifo_inst/buff[115][2] ), .I1(\i11/fifo_inst/buff[113][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3499.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3500 (.I0(n2044), .I1(n2043), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1785), .O(n2045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3500.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3501 (.I0(n2042), .I1(n2041), .I2(n2045), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__3501.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__3502 (.I0(\i11/fifo_inst/buff[123][2] ), .I1(\i11/fifo_inst/buff[121][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3502.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3503 (.I0(\i11/fifo_inst/buff[120][2] ), .I1(\i11/fifo_inst/buff[122][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3503.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3504 (.I0(\i11/fifo_inst/buff[124][2] ), .I1(\i11/fifo_inst/buff[126][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3504.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3505 (.I0(\i11/fifo_inst/buff[127][2] ), .I1(\i11/fifo_inst/buff[125][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2049), .O(n2050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3505.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3506 (.I0(n2048), .I1(n2047), .I2(n2050), .I3(n1785), 
            .O(n2051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3506.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3507 (.I0(n2051), .I1(n2046), .I2(n1795), .I3(n1829), 
            .O(n2052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3507.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3508 (.I0(\i11/fifo_inst/buff[76][2] ), .I1(\i11/fifo_inst/buff[78][2] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__3508.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__3509 (.I0(\i11/fifo_inst/buff[79][2] ), .I1(\i11/fifo_inst/buff[77][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n2054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__3509.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__3510 (.I0(\i11/fifo_inst/buff[72][2] ), .I1(\i11/fifo_inst/buff[74][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3510.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3511 (.I0(\i11/fifo_inst/buff[75][2] ), .I1(\i11/fifo_inst/buff[73][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3511.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3512 (.I0(n2056), .I1(n2055), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1785), .O(n2057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3512.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3513 (.I0(n2054), .I1(n2053), .I2(n2057), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__3513.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__3514 (.I0(\i11/fifo_inst/buff[67][2] ), .I1(\i11/fifo_inst/buff[65][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3514.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3515 (.I0(\i11/fifo_inst/buff[64][2] ), .I1(\i11/fifo_inst/buff[66][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3515.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3516 (.I0(\i11/fifo_inst/buff[68][2] ), .I1(\i11/fifo_inst/buff[70][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3516.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3517 (.I0(\i11/fifo_inst/buff[71][2] ), .I1(\i11/fifo_inst/buff[69][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2061), .O(n2062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3517.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3518 (.I0(n2060), .I1(n2059), .I2(n2062), .I3(n1785), 
            .O(n2063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3518.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3519 (.I0(n2063), .I1(n2058), .I2(n1822), .I3(n1795), 
            .O(n2064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3519.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3520 (.I0(\i11/fifo_inst/buff[92][2] ), .I1(\i11/fifo_inst/buff[94][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3520.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3521 (.I0(\i11/fifo_inst/buff[93][2] ), .I1(\i11/fifo_inst/buff[95][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2065), .O(n2066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__3521.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__3522 (.I0(\i11/fifo_inst/buff[88][2] ), .I1(\i11/fifo_inst/buff[90][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3522.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3523 (.I0(\i11/fifo_inst/buff[91][2] ), .I1(\i11/fifo_inst/buff[89][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2067), .O(n2068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3523.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3524 (.I0(n2068), .I1(n2066), .I2(n1795), .I3(n1785), 
            .O(n2069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__3524.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__3525 (.I0(\i11/fifo_inst/buff[80][2] ), .I1(\i11/fifo_inst/buff[82][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3525.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3526 (.I0(\i11/fifo_inst/buff[83][2] ), .I1(\i11/fifo_inst/buff[81][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3526.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3527 (.I0(n2071), .I1(n2070), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1785), .O(n2072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3527.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3528 (.I0(\i11/fifo_inst/buff[86][2] ), .I1(\i11/fifo_inst/buff[84][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n2073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__3528.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__3529 (.I0(\i11/fifo_inst/buff[87][2] ), .I1(\i11/fifo_inst/buff[85][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3529.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3530 (.I0(n2074), .I1(n1819), .I2(n2073), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__3530.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__3531 (.I0(n2072), .I1(n2075), .I2(n1795), .I3(n1808), 
            .O(n2076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__3531.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__3532 (.I0(\i11/fifo_inst/buff[96][2] ), .I1(\i11/fifo_inst/buff[98][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3532.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3533 (.I0(\i11/fifo_inst/buff[99][2] ), .I1(\i11/fifo_inst/buff[97][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3533.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3534 (.I0(n2078), .I1(n2077), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1785), .O(n2079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3534.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3535 (.I0(\i11/fifo_inst/buff[102][2] ), .I1(\i11/fifo_inst/buff[100][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n2080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__3535.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__3536 (.I0(\i11/fifo_inst/buff[103][2] ), .I1(\i11/fifo_inst/buff[101][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3536.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3537 (.I0(n2081), .I1(n1819), .I2(n2080), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__3537.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__3538 (.I0(n2079), .I1(n2082), .I2(n1795), .I3(n1794), 
            .O(n2083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__3538.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__3539 (.I0(\i11/fifo_inst/buff[108][2] ), .I1(\i11/fifo_inst/buff[110][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3539.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3540 (.I0(\i11/fifo_inst/buff[109][2] ), .I1(\i11/fifo_inst/buff[111][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2084), .O(n2085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__3540.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__3541 (.I0(\i11/fifo_inst/buff[104][2] ), .I1(\i11/fifo_inst/buff[106][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3541.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3542 (.I0(\i11/fifo_inst/buff[107][2] ), .I1(\i11/fifo_inst/buff[105][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2086), .O(n2087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3542.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3543 (.I0(n2087), .I1(n2085), .I2(n1795), .I3(n1785), 
            .O(n2088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__3543.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__3544 (.I0(n2088), .I1(n2083), .I2(n2069), .I3(n2076), 
            .O(n2089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__3544.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__3545 (.I0(n2064), .I1(n2052), .I2(n2089), .I3(n1895), 
            .O(n2090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__3545.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__3546 (.I0(n1780), .I1(\rx_d[2] ), .O(n2091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3546.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3547 (.I0(n2040), .I1(n1838), .I2(n2090), .I3(n2091), 
            .O(\fifo_inst/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4 */ ;
    defparam LUT__3547.LUTMASK = 16'hfff4;
    EFX_LUT4 LUT__3548 (.I0(\i11/fifo_inst/buff[67][3] ), .I1(\i11/fifo_inst/buff[65][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3548.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3549 (.I0(\i11/fifo_inst/buff[64][3] ), .I1(\i11/fifo_inst/buff[66][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3549.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3550 (.I0(\i11/fifo_inst/buff[68][3] ), .I1(\i11/fifo_inst/buff[70][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3550.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3551 (.I0(\i11/fifo_inst/buff[71][3] ), .I1(\i11/fifo_inst/buff[69][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2094), .O(n2095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3551.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3552 (.I0(n2093), .I1(n2092), .I2(n2095), .I3(n1785), 
            .O(n2096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3552.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3553 (.I0(\i11/fifo_inst/buff[75][3] ), .I1(\i11/fifo_inst/buff[73][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3553.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3554 (.I0(\i11/fifo_inst/buff[72][3] ), .I1(\i11/fifo_inst/buff[74][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3554.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3555 (.I0(\i11/fifo_inst/buff[76][3] ), .I1(\i11/fifo_inst/buff[78][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3555.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3556 (.I0(\i11/fifo_inst/buff[79][3] ), .I1(\i11/fifo_inst/buff[77][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2099), .O(n2100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3556.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3557 (.I0(n2098), .I1(n2097), .I2(n2100), .I3(n1785), 
            .O(n2101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3557.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3558 (.I0(n2101), .I1(n2096), .I2(n1822), .I3(n1795), 
            .O(n2102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3558.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3559 (.I0(\i11/fifo_inst/buff[116][3] ), .I1(\i11/fifo_inst/buff[118][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3559.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3560 (.I0(\i11/fifo_inst/buff[119][3] ), .I1(\i11/fifo_inst/buff[117][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3560.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3561 (.I0(\i11/fifo_inst/buff[112][3] ), .I1(\i11/fifo_inst/buff[114][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3561.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3562 (.I0(\i11/fifo_inst/buff[115][3] ), .I1(\i11/fifo_inst/buff[113][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2105), .O(n2106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3562.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3563 (.I0(n2104), .I1(n2103), .I2(n2106), .I3(n1785), 
            .O(n2107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3563.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3564 (.I0(\i11/fifo_inst/buff[123][3] ), .I1(\i11/fifo_inst/buff[121][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3564.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3565 (.I0(\i11/fifo_inst/buff[120][3] ), .I1(\i11/fifo_inst/buff[122][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3565.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3566 (.I0(\i11/fifo_inst/buff[124][3] ), .I1(\i11/fifo_inst/buff[126][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3566.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3567 (.I0(\i11/fifo_inst/buff[127][3] ), .I1(\i11/fifo_inst/buff[125][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2110), .O(n2111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3567.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3568 (.I0(n2109), .I1(n2108), .I2(n2111), .I3(n1785), 
            .O(n2112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3568.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3569 (.I0(n2112), .I1(n2107), .I2(n1795), .I3(n1829), 
            .O(n2113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3569.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3570 (.I0(\i11/fifo_inst/buff[100][3] ), .I1(\i11/fifo_inst/buff[102][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3570.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3571 (.I0(\i11/fifo_inst/buff[103][3] ), .I1(\i11/fifo_inst/buff[101][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2114), .O(n2115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3571.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3572 (.I0(\i11/fifo_inst/buff[96][3] ), .I1(\i11/fifo_inst/buff[98][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3572.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3573 (.I0(\i11/fifo_inst/buff[99][3] ), .I1(\i11/fifo_inst/buff[97][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2116), .O(n2117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3573.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3574 (.I0(n2117), .I1(n2115), .I2(n1785), .I3(n1795), 
            .O(n2118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3574.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3575 (.I0(\i11/fifo_inst/buff[111][3] ), .I1(\i11/fifo_inst/buff[109][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n2119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__3575.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__3576 (.I0(\i11/fifo_inst/buff[108][3] ), .I1(\i11/fifo_inst/buff[110][3] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__3576.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__3577 (.I0(n2119), .I1(n2120), .I2(n1795), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__3577.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__3578 (.I0(\i11/fifo_inst/buff[104][3] ), .I1(\i11/fifo_inst/buff[106][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3578.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3579 (.I0(\i11/fifo_inst/buff[107][3] ), .I1(\i11/fifo_inst/buff[105][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2122), .O(n2123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3579.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3580 (.I0(n2123), .I1(n1785), .I2(n2121), .I3(n1794), 
            .O(n2124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__3580.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__3581 (.I0(\i11/fifo_inst/buff[84][3] ), .I1(\i11/fifo_inst/buff[86][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3581.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3582 (.I0(\i11/fifo_inst/buff[87][3] ), .I1(\i11/fifo_inst/buff[85][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2125), .O(n2126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3582.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3583 (.I0(\i11/fifo_inst/buff[80][3] ), .I1(\i11/fifo_inst/buff[82][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3583.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3584 (.I0(\i11/fifo_inst/buff[83][3] ), .I1(\i11/fifo_inst/buff[81][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2127), .O(n2128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3584.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3585 (.I0(n2128), .I1(n2126), .I2(n1785), .I3(n1795), 
            .O(n2129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3585.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3586 (.I0(\i11/fifo_inst/buff[95][3] ), .I1(\i11/fifo_inst/buff[93][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n2130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__3586.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__3587 (.I0(\i11/fifo_inst/buff[92][3] ), .I1(\i11/fifo_inst/buff[94][3] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__3587.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__3588 (.I0(n2130), .I1(n2131), .I2(n1795), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__3588.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__3589 (.I0(\i11/fifo_inst/buff[88][3] ), .I1(\i11/fifo_inst/buff[90][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3589.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3590 (.I0(\i11/fifo_inst/buff[91][3] ), .I1(\i11/fifo_inst/buff[89][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2133), .O(n2134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3590.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3591 (.I0(n2134), .I1(n1785), .I2(n2132), .I3(n1808), 
            .O(n2135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__3591.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__3592 (.I0(n2129), .I1(n2135), .I2(n2118), .I3(n2124), 
            .O(n2136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__3592.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__3593 (.I0(n2102), .I1(n2113), .I2(n2136), .I3(n1895), 
            .O(n2137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__3593.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__3594 (.I0(rx_en_fifo), .I1(n1745), .I2(\rx_d[3] ), .O(n2138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3594.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3595 (.I0(\i11/fifo_inst/buff[40][3] ), .I1(\i11/fifo_inst/buff[42][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3595.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3596 (.I0(\i11/fifo_inst/buff[43][3] ), .I1(\i11/fifo_inst/buff[41][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2139), .O(n2140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3596.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3597 (.I0(\i11/fifo_inst/buff[44][3] ), .I1(\i11/fifo_inst/buff[46][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3597.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3598 (.I0(\i11/fifo_inst/buff[47][3] ), .I1(\i11/fifo_inst/buff[45][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2141), .O(n2142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3598.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3599 (.I0(\i11/fifo_inst/buff[36][3] ), .I1(\i11/fifo_inst/buff[38][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3599.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3600 (.I0(\i11/fifo_inst/buff[39][3] ), .I1(\i11/fifo_inst/buff[37][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3600.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3601 (.I0(n2144), .I1(n2143), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n2145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3601.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3602 (.I0(\i11/fifo_inst/buff[32][3] ), .I1(\i11/fifo_inst/buff[34][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3602.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3603 (.I0(\i11/fifo_inst/buff[35][3] ), .I1(\i11/fifo_inst/buff[33][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3603.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3604 (.I0(n2147), .I1(n2146), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3604.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3605 (.I0(n1853), .I1(n2142), .I2(n2145), .I3(n2148), 
            .O(n2149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__3605.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__3606 (.I0(n1865), .I1(n2140), .I2(n2149), .I3(n1794), 
            .O(n2150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__3606.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__3607 (.I0(\i11/fifo_inst/buff[51][3] ), .I1(\i11/fifo_inst/buff[49][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3607.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3608 (.I0(\i11/fifo_inst/buff[48][3] ), .I1(\i11/fifo_inst/buff[50][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3608.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3609 (.I0(\i11/fifo_inst/buff[52][3] ), .I1(\i11/fifo_inst/buff[54][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3609.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3610 (.I0(\i11/fifo_inst/buff[55][3] ), .I1(\i11/fifo_inst/buff[53][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2153), .O(n2154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3610.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3611 (.I0(n2152), .I1(n2151), .I2(n2154), .I3(n1785), 
            .O(n2155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3611.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3612 (.I0(\i11/fifo_inst/buff[59][3] ), .I1(\i11/fifo_inst/buff[57][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3612.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3613 (.I0(\i11/fifo_inst/buff[56][3] ), .I1(\i11/fifo_inst/buff[58][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3613.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3614 (.I0(\i11/fifo_inst/buff[60][3] ), .I1(\i11/fifo_inst/buff[62][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3614.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3615 (.I0(\i11/fifo_inst/buff[63][3] ), .I1(\i11/fifo_inst/buff[61][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2158), .O(n2159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3615.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3616 (.I0(n2157), .I1(n2156), .I2(n2159), .I3(n1785), 
            .O(n2160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3616.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3617 (.I0(n2160), .I1(n2155), .I2(n1795), .I3(n1829), 
            .O(n2161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3617.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3618 (.I0(\i11/fifo_inst/buff[11][3] ), .I1(\i11/fifo_inst/buff[9][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3618.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3619 (.I0(\i11/fifo_inst/buff[8][3] ), .I1(\i11/fifo_inst/buff[10][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3619.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3620 (.I0(\i11/fifo_inst/buff[24][3] ), .I1(\i11/fifo_inst/buff[26][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3620.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3621 (.I0(\i11/fifo_inst/buff[27][3] ), .I1(\i11/fifo_inst/buff[25][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2164), .O(n2165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3621.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3622 (.I0(n2163), .I1(n2162), .I2(n2165), .I3(n1882), 
            .O(n2166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3622.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3623 (.I0(\i11/fifo_inst/buff[0][3] ), .I1(\i11/fifo_inst/buff[2][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3623.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3624 (.I0(\i11/fifo_inst/buff[3][3] ), .I1(\i11/fifo_inst/buff[1][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2167), .O(n2168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3624.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3625 (.I0(\i11/fifo_inst/buff[16][3] ), .I1(\i11/fifo_inst/buff[18][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3625.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3626 (.I0(\i11/fifo_inst/buff[19][3] ), .I1(\i11/fifo_inst/buff[17][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2169), .O(n2170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3626.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3627 (.I0(n2170), .I1(n2168), .I2(n1882), .I3(n1795), 
            .O(n2171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3627.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3628 (.I0(n1795), .I1(n2166), .I2(n2171), .I3(n1785), 
            .O(n2172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__3628.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__3629 (.I0(\i11/fifo_inst/buff[15][3] ), .I1(\i11/fifo_inst/buff[13][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3629.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3630 (.I0(\i11/fifo_inst/buff[12][3] ), .I1(\i11/fifo_inst/buff[14][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3630.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3631 (.I0(\i11/fifo_inst/buff[28][3] ), .I1(\i11/fifo_inst/buff[30][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3631.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3632 (.I0(\i11/fifo_inst/buff[31][3] ), .I1(\i11/fifo_inst/buff[29][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2175), .O(n2176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3632.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3633 (.I0(n2174), .I1(n2173), .I2(n2176), .I3(n1882), 
            .O(n2177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3633.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3634 (.I0(\i11/fifo_inst/buff[4][3] ), .I1(\i11/fifo_inst/buff[6][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3634.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3635 (.I0(\i11/fifo_inst/buff[7][3] ), .I1(\i11/fifo_inst/buff[5][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2178), .O(n2179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3635.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3636 (.I0(\i11/fifo_inst/buff[20][3] ), .I1(\i11/fifo_inst/buff[22][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3636.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3637 (.I0(\i11/fifo_inst/buff[23][3] ), .I1(\i11/fifo_inst/buff[21][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2180), .O(n2181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3637.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3638 (.I0(n2181), .I1(n2179), .I2(n1882), .I3(n1861), 
            .O(n2182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3638.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3639 (.I0(n2177), .I1(n1853), .I2(n2182), .I3(n1881), 
            .O(n2183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__3639.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__3640 (.I0(n2183), .I1(n2172), .I2(n2150), .I3(n2161), 
            .O(n2184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__3640.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__3641 (.I0(n2184), .I1(n1838), .I2(n2138), .I3(n2137), 
            .O(\fifo_inst/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4 */ ;
    defparam LUT__3641.LUTMASK = 16'hfff4;
    EFX_LUT4 LUT__3642 (.I0(\i11/fifo_inst/buff[84][4] ), .I1(\i11/fifo_inst/buff[86][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3642.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3643 (.I0(\i11/fifo_inst/buff[87][4] ), .I1(\i11/fifo_inst/buff[85][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2185), .O(n2186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3643.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3644 (.I0(\i11/fifo_inst/buff[116][4] ), .I1(\i11/fifo_inst/buff[118][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3644.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3645 (.I0(\i11/fifo_inst/buff[119][4] ), .I1(\i11/fifo_inst/buff[117][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2187), .O(n2188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3645.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3646 (.I0(n2188), .I1(n2186), .I2(n1785), .I3(n1881), 
            .O(n2189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3646.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3647 (.I0(\i11/fifo_inst/buff[80][4] ), .I1(\i11/fifo_inst/buff[82][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3647.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3648 (.I0(\i11/fifo_inst/buff[83][4] ), .I1(\i11/fifo_inst/buff[81][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2190), .O(n2191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3648.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3649 (.I0(\i11/fifo_inst/buff[112][4] ), .I1(\i11/fifo_inst/buff[114][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3649.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3650 (.I0(\i11/fifo_inst/buff[115][4] ), .I1(\i11/fifo_inst/buff[113][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2192), .O(n2193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3650.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3651 (.I0(n2193), .I1(n2191), .I2(n1881), .I3(n1785), 
            .O(n2194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3651.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3652 (.I0(n2189), .I1(n2194), .I2(n1795), .O(n2195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3652.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3653 (.I0(\i11/fifo_inst/buff[92][4] ), .I1(\i11/fifo_inst/buff[94][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3653.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3654 (.I0(\i11/fifo_inst/buff[95][4] ), .I1(\i11/fifo_inst/buff[93][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2196), .O(n2197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3654.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3655 (.I0(\i11/fifo_inst/buff[124][4] ), .I1(\i11/fifo_inst/buff[126][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3655.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3656 (.I0(\i11/fifo_inst/buff[127][4] ), .I1(\i11/fifo_inst/buff[125][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2198), .O(n2199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3656.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3657 (.I0(n2199), .I1(n2197), .I2(n1785), .I3(n1881), 
            .O(n2200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3657.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3658 (.I0(\i11/fifo_inst/buff[88][4] ), .I1(\i11/fifo_inst/buff[90][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3658.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3659 (.I0(\i11/fifo_inst/buff[91][4] ), .I1(\i11/fifo_inst/buff[89][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2201), .O(n2202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3659.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3660 (.I0(\i11/fifo_inst/buff[120][4] ), .I1(\i11/fifo_inst/buff[122][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3660.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3661 (.I0(\i11/fifo_inst/buff[123][4] ), .I1(\i11/fifo_inst/buff[121][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2203), .O(n2204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3661.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3662 (.I0(n2204), .I1(n2202), .I2(n1881), .I3(n1785), 
            .O(n2205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3662.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3663 (.I0(n2200), .I1(n2205), .I2(n1795), .O(n2206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__3663.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__3664 (.I0(\i11/fifo_inst/buff[64][4] ), .I1(\i11/fifo_inst/buff[66][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3664.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3665 (.I0(\i11/fifo_inst/buff[67][4] ), .I1(\i11/fifo_inst/buff[65][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3665.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3666 (.I0(n2208), .I1(n2207), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3666.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3667 (.I0(\i11/fifo_inst/buff[76][4] ), .I1(\i11/fifo_inst/buff[78][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3667.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3668 (.I0(\i11/fifo_inst/buff[79][4] ), .I1(\i11/fifo_inst/buff[77][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3668.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3669 (.I0(n2211), .I1(n2210), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1853), .O(n2212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3669.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3670 (.I0(\i11/fifo_inst/buff[68][4] ), .I1(\i11/fifo_inst/buff[70][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3670.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3671 (.I0(\i11/fifo_inst/buff[71][4] ), .I1(\i11/fifo_inst/buff[69][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3671.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3672 (.I0(n2214), .I1(n2213), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n2215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3672.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3673 (.I0(\i11/fifo_inst/buff[72][4] ), .I1(\i11/fifo_inst/buff[74][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3673.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3674 (.I0(\i11/fifo_inst/buff[75][4] ), .I1(\i11/fifo_inst/buff[73][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3674.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3675 (.I0(n2217), .I1(n2216), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3675.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3676 (.I0(n2209), .I1(n2212), .I2(n2215), .I3(n2218), 
            .O(n2219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3676.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3677 (.I0(\i11/fifo_inst/buff[100][4] ), .I1(\i11/fifo_inst/buff[102][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3677.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3678 (.I0(\i11/fifo_inst/buff[103][4] ), .I1(\i11/fifo_inst/buff[101][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3678.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3679 (.I0(n2221), .I1(n2220), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n2222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3679.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3680 (.I0(\i11/fifo_inst/buff[108][4] ), .I1(\i11/fifo_inst/buff[110][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3680.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3681 (.I0(\i11/fifo_inst/buff[111][4] ), .I1(\i11/fifo_inst/buff[109][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3681.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3682 (.I0(n2224), .I1(n2223), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1853), .O(n2225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3682.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3683 (.I0(\i11/fifo_inst/buff[96][4] ), .I1(\i11/fifo_inst/buff[98][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3683.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3684 (.I0(\i11/fifo_inst/buff[99][4] ), .I1(\i11/fifo_inst/buff[97][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3684.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3685 (.I0(n2227), .I1(n2226), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3685.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3686 (.I0(\i11/fifo_inst/buff[104][4] ), .I1(\i11/fifo_inst/buff[106][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3686.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3687 (.I0(\i11/fifo_inst/buff[107][4] ), .I1(\i11/fifo_inst/buff[105][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3687.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3688 (.I0(n2230), .I1(n2229), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3688.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3689 (.I0(n2222), .I1(n2225), .I2(n2228), .I3(n2231), 
            .O(n2232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3689.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3690 (.I0(n2232), .I1(n2219), .I2(n1881), .O(n2233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3690.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3691 (.I0(n2206), .I1(n2195), .I2(n2233), .I3(n1882), 
            .O(n2234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3691.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3692 (.I0(n1780), .I1(\rx_d[4] ), .O(n2235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3692.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3693 (.I0(\i11/fifo_inst/buff[4][4] ), .I1(\i11/fifo_inst/buff[6][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3693.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3694 (.I0(\i11/fifo_inst/buff[7][4] ), .I1(\i11/fifo_inst/buff[5][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2236), .O(n2237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3694.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3695 (.I0(\i11/fifo_inst/buff[20][4] ), .I1(\i11/fifo_inst/buff[22][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3695.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3696 (.I0(\i11/fifo_inst/buff[23][4] ), .I1(\i11/fifo_inst/buff[21][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2238), .O(n2239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3696.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3697 (.I0(n2239), .I1(n2237), .I2(n1882), .I3(n1861), 
            .O(n2240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3697.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3698 (.I0(\i11/fifo_inst/buff[8][4] ), .I1(\i11/fifo_inst/buff[10][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3698.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3699 (.I0(\i11/fifo_inst/buff[11][4] ), .I1(\i11/fifo_inst/buff[9][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2241), .O(n2242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3699.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3700 (.I0(\i11/fifo_inst/buff[24][4] ), .I1(\i11/fifo_inst/buff[26][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3700.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3701 (.I0(\i11/fifo_inst/buff[27][4] ), .I1(\i11/fifo_inst/buff[25][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2243), .O(n2244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3701.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3702 (.I0(n2244), .I1(n2242), .I2(n1865), .I3(n1882), 
            .O(n2245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3702.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3703 (.I0(n1778), .I1(n1837), .I2(n1881), .I3(ceg_net146), 
            .O(n2246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__3703.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__3704 (.I0(n2240), .I1(n2245), .I2(n2246), .O(n2247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3704.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3705 (.I0(\i11/fifo_inst/buff[12][4] ), .I1(\i11/fifo_inst/buff[14][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3705.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3706 (.I0(\i11/fifo_inst/buff[15][4] ), .I1(\i11/fifo_inst/buff[13][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2248), .O(n2249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3706.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3707 (.I0(\i11/fifo_inst/buff[28][4] ), .I1(\i11/fifo_inst/buff[30][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3707.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3708 (.I0(\i11/fifo_inst/buff[31][4] ), .I1(\i11/fifo_inst/buff[29][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2250), .O(n2251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3708.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3709 (.I0(n2251), .I1(n2249), .I2(n1882), .O(n2252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3709.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3710 (.I0(\i11/fifo_inst/buff[0][4] ), .I1(\i11/fifo_inst/buff[2][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3710.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3711 (.I0(\i11/fifo_inst/buff[3][4] ), .I1(\i11/fifo_inst/buff[1][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2253), .O(n2254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3711.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3712 (.I0(\i11/fifo_inst/buff[16][4] ), .I1(\i11/fifo_inst/buff[18][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3712.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3713 (.I0(\i11/fifo_inst/buff[19][4] ), .I1(\i11/fifo_inst/buff[17][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2255), .O(n2256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3713.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3714 (.I0(n2256), .I1(n2254), .I2(n1882), .O(n2257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3714.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3715 (.I0(n1857), .I1(n2257), .I2(n2252), .I3(n1853), 
            .O(n2258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__3715.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__3716 (.I0(\i11/fifo_inst/buff[56][4] ), .I1(\i11/fifo_inst/buff[58][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3716.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3717 (.I0(\i11/fifo_inst/buff[59][4] ), .I1(\i11/fifo_inst/buff[57][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3717.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3718 (.I0(n2260), .I1(n2259), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3718.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3719 (.I0(\i11/fifo_inst/buff[60][4] ), .I1(\i11/fifo_inst/buff[62][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3719.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3720 (.I0(\i11/fifo_inst/buff[63][4] ), .I1(\i11/fifo_inst/buff[61][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3720.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3721 (.I0(n2263), .I1(n2262), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1853), .O(n2264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3721.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3722 (.I0(\i11/fifo_inst/buff[48][4] ), .I1(\i11/fifo_inst/buff[50][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3722.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3723 (.I0(\i11/fifo_inst/buff[51][4] ), .I1(\i11/fifo_inst/buff[49][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3723.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3724 (.I0(n2266), .I1(n2265), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3724.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3725 (.I0(\i11/fifo_inst/buff[52][4] ), .I1(\i11/fifo_inst/buff[54][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3725.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3726 (.I0(\i11/fifo_inst/buff[55][4] ), .I1(\i11/fifo_inst/buff[53][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3726.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3727 (.I0(n2269), .I1(n2268), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n2270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3727.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3728 (.I0(n2261), .I1(n2264), .I2(n2267), .I3(n2270), 
            .O(n2271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3728.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3729 (.I0(n2271), .I1(n1838), .I2(n1829), .O(n2272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3729.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3730 (.I0(\i11/fifo_inst/buff[44][4] ), .I1(\i11/fifo_inst/buff[46][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3730.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3731 (.I0(\i11/fifo_inst/buff[47][4] ), .I1(\i11/fifo_inst/buff[45][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2273), .O(n2274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3731.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3732 (.I0(\i11/fifo_inst/buff[36][4] ), .I1(\i11/fifo_inst/buff[38][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3732.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3733 (.I0(\i11/fifo_inst/buff[39][4] ), .I1(\i11/fifo_inst/buff[37][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2275), .O(n2276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3733.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3734 (.I0(n2276), .I1(n2274), .I2(n1785), .I3(n1795), 
            .O(n2277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3734.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3735 (.I0(\i11/fifo_inst/buff[40][4] ), .I1(\i11/fifo_inst/buff[42][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3735.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3736 (.I0(\i11/fifo_inst/buff[43][4] ), .I1(\i11/fifo_inst/buff[41][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2278), .O(n2279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3736.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3737 (.I0(\i11/fifo_inst/buff[32][4] ), .I1(\i11/fifo_inst/buff[34][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3737.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3738 (.I0(\i11/fifo_inst/buff[35][4] ), .I1(\i11/fifo_inst/buff[33][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2280), .O(n2281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3738.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3739 (.I0(n2281), .I1(n2279), .I2(n1795), .I3(n1785), 
            .O(n2282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3739.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3740 (.I0(n2277), .I1(n2282), .I2(n1794), .I3(n1838), 
            .O(n2283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3740.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3741 (.I0(n2258), .I1(n2247), .I2(n2272), .I3(n2283), 
            .O(n2284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__3741.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__3742 (.I0(n2234), .I1(n1895), .I2(n2235), .I3(n2284), 
            .O(\fifo_inst/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8ff */ ;
    defparam LUT__3742.LUTMASK = 16'hf8ff;
    EFX_LUT4 LUT__3743 (.I0(\i11/fifo_inst/buff[64][5] ), .I1(\i11/fifo_inst/buff[66][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3743.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3744 (.I0(\i11/fifo_inst/buff[67][5] ), .I1(\i11/fifo_inst/buff[65][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2285), .O(n2286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3744.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3745 (.I0(\i11/fifo_inst/buff[72][5] ), .I1(\i11/fifo_inst/buff[74][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3745.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3746 (.I0(\i11/fifo_inst/buff[75][5] ), .I1(\i11/fifo_inst/buff[73][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2287), .O(n2288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3746.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3747 (.I0(\i11/fifo_inst/buff[76][5] ), .I1(\i11/fifo_inst/buff[78][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3747.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3748 (.I0(\i11/fifo_inst/buff[79][5] ), .I1(\i11/fifo_inst/buff[77][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3748.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3749 (.I0(n2290), .I1(n2289), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1853), .O(n2291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3749.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3750 (.I0(\i11/fifo_inst/buff[68][5] ), .I1(\i11/fifo_inst/buff[70][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3750.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3751 (.I0(\i11/fifo_inst/buff[71][5] ), .I1(\i11/fifo_inst/buff[69][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3751.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3752 (.I0(n2293), .I1(n2292), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n2294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3752.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3753 (.I0(n1865), .I1(n2288), .I2(n2291), .I3(n2294), 
            .O(n2295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__3753.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__3754 (.I0(n1857), .I1(n2286), .I2(n2295), .I3(n1822), 
            .O(n2296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__3754.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__3755 (.I0(\i11/fifo_inst/buff[103][5] ), .I1(\i11/fifo_inst/buff[101][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3755.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3756 (.I0(\i11/fifo_inst/buff[100][5] ), .I1(\i11/fifo_inst/buff[102][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3756.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3757 (.I0(\i11/fifo_inst/buff[96][5] ), .I1(\i11/fifo_inst/buff[98][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3757.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3758 (.I0(\i11/fifo_inst/buff[99][5] ), .I1(\i11/fifo_inst/buff[97][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2299), .O(n2300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3758.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3759 (.I0(n2298), .I1(n2297), .I2(n2300), .I3(n1785), 
            .O(n2301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__3759.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__3760 (.I0(\i11/fifo_inst/buff[111][5] ), .I1(\i11/fifo_inst/buff[109][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3760.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3761 (.I0(\i11/fifo_inst/buff[108][5] ), .I1(\i11/fifo_inst/buff[110][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3761.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3762 (.I0(\i11/fifo_inst/buff[104][5] ), .I1(\i11/fifo_inst/buff[106][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3762.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3763 (.I0(\i11/fifo_inst/buff[107][5] ), .I1(\i11/fifo_inst/buff[105][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2304), .O(n2305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3763.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3764 (.I0(n2303), .I1(n2302), .I2(n2305), .I3(n1785), 
            .O(n2306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__3764.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__3765 (.I0(n2306), .I1(n2301), .I2(n1794), .I3(n1795), 
            .O(n2307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3765.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3766 (.I0(\i11/fifo_inst/buff[95][5] ), .I1(\i11/fifo_inst/buff[93][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3766.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3767 (.I0(\i11/fifo_inst/buff[92][5] ), .I1(\i11/fifo_inst/buff[94][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3767.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3768 (.I0(\i11/fifo_inst/buff[124][5] ), .I1(\i11/fifo_inst/buff[126][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3768.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3769 (.I0(\i11/fifo_inst/buff[127][5] ), .I1(\i11/fifo_inst/buff[125][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2310), .O(n2311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3769.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3770 (.I0(n2309), .I1(n2308), .I2(n2311), .I3(n1881), 
            .O(n2312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3770.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3771 (.I0(\i11/fifo_inst/buff[91][5] ), .I1(\i11/fifo_inst/buff[89][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3771.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3772 (.I0(\i11/fifo_inst/buff[88][5] ), .I1(\i11/fifo_inst/buff[90][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3772.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3773 (.I0(\i11/fifo_inst/buff[120][5] ), .I1(\i11/fifo_inst/buff[122][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3773.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3774 (.I0(\i11/fifo_inst/buff[123][5] ), .I1(\i11/fifo_inst/buff[121][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2315), .O(n2316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3774.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3775 (.I0(n2314), .I1(n2313), .I2(n2316), .I3(n1881), 
            .O(n2317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3775.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3776 (.I0(n2317), .I1(n2312), .I2(n1795), .I3(n1785), 
            .O(n2318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__3776.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__3777 (.I0(\i11/fifo_inst/buff[87][5] ), .I1(\i11/fifo_inst/buff[85][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3777.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3778 (.I0(\i11/fifo_inst/buff[84][5] ), .I1(\i11/fifo_inst/buff[86][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3778.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3779 (.I0(\i11/fifo_inst/buff[83][5] ), .I1(\i11/fifo_inst/buff[81][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3779.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3780 (.I0(\i11/fifo_inst/buff[80][5] ), .I1(\i11/fifo_inst/buff[82][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3780.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3781 (.I0(n2322), .I1(n2321), .I2(n1785), .I3(\fifo_inst/rd_index[5] ), 
            .O(n2323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__3781.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__3782 (.I0(n2320), .I1(n1785), .I2(n2319), .I3(n2323), 
            .O(n2324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__3782.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__3783 (.I0(\i11/fifo_inst/buff[116][5] ), .I1(\i11/fifo_inst/buff[118][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3783.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3784 (.I0(\i11/fifo_inst/buff[119][5] ), .I1(\i11/fifo_inst/buff[117][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2325), .O(n2326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3784.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3785 (.I0(\i11/fifo_inst/buff[112][5] ), .I1(\i11/fifo_inst/buff[114][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3785.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3786 (.I0(\i11/fifo_inst/buff[115][5] ), .I1(\i11/fifo_inst/buff[113][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2327), .O(n2328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3786.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3787 (.I0(n2328), .I1(n2326), .I2(n1785), .I3(\fifo_inst/rd_index[5] ), 
            .O(n2329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3787.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3788 (.I0(n2329), .I1(n2324), .I2(n1795), .I3(n1882), 
            .O(n2330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__3788.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__3789 (.I0(n2330), .I1(n2318), .I2(n2296), .I3(n2307), 
            .O(n2331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__3789.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__3790 (.I0(\i11/fifo_inst/buff[47][5] ), .I1(\i11/fifo_inst/buff[45][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3790.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3791 (.I0(\i11/fifo_inst/buff[44][5] ), .I1(\i11/fifo_inst/buff[46][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3791.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3792 (.I0(\i11/fifo_inst/buff[60][5] ), .I1(\i11/fifo_inst/buff[62][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3792.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3793 (.I0(\i11/fifo_inst/buff[63][5] ), .I1(\i11/fifo_inst/buff[61][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2334), .O(n2335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3793.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3794 (.I0(n2333), .I1(n2332), .I2(n2335), .I3(n1882), 
            .O(n2336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3794.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3795 (.I0(\i11/fifo_inst/buff[43][5] ), .I1(\i11/fifo_inst/buff[41][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3795.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3796 (.I0(\i11/fifo_inst/buff[40][5] ), .I1(\i11/fifo_inst/buff[42][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3796.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3797 (.I0(\i11/fifo_inst/buff[56][5] ), .I1(\i11/fifo_inst/buff[58][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3797.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3798 (.I0(\i11/fifo_inst/buff[59][5] ), .I1(\i11/fifo_inst/buff[57][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2339), .O(n2340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3798.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3799 (.I0(n2338), .I1(n2337), .I2(n2340), .I3(n1882), 
            .O(n2341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3799.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3800 (.I0(n2341), .I1(n2336), .I2(n1795), .I3(n1785), 
            .O(n2342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3800.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3801 (.I0(\i11/fifo_inst/buff[39][5] ), .I1(\i11/fifo_inst/buff[37][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3801.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3802 (.I0(\i11/fifo_inst/buff[36][5] ), .I1(\i11/fifo_inst/buff[38][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3802.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3803 (.I0(\i11/fifo_inst/buff[52][5] ), .I1(\i11/fifo_inst/buff[54][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3803.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3804 (.I0(\i11/fifo_inst/buff[55][5] ), .I1(\i11/fifo_inst/buff[53][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2345), .O(n2346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3804.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3805 (.I0(n2344), .I1(n2343), .I2(n2346), .I3(n1882), 
            .O(n2347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__3805.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__3806 (.I0(\i11/fifo_inst/buff[32][5] ), .I1(\i11/fifo_inst/buff[34][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3806.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3807 (.I0(\i11/fifo_inst/buff[35][5] ), .I1(\i11/fifo_inst/buff[33][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2348), .O(n2349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3807.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3808 (.I0(\i11/fifo_inst/buff[48][5] ), .I1(\i11/fifo_inst/buff[50][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3808.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3809 (.I0(\i11/fifo_inst/buff[51][5] ), .I1(\i11/fifo_inst/buff[49][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2350), .O(n2351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3809.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3810 (.I0(n2351), .I1(n2349), .I2(n1882), .I3(n1785), 
            .O(n2352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3810.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3811 (.I0(n2347), .I1(n1785), .I2(n2352), .I3(n1795), 
            .O(n2353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__3811.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__3812 (.I0(n2353), .I1(n2342), .I2(n1881), .I3(n1838), 
            .O(n2354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__3812.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__3813 (.I0(\i11/fifo_inst/buff[2][5] ), .I1(\i11/fifo_inst/buff[0][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3813.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3814 (.I0(\i11/fifo_inst/buff[1][5] ), .I1(\i11/fifo_inst/buff[3][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3814.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3815 (.I0(n2356), .I1(n2355), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3815.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3816 (.I0(\i11/fifo_inst/buff[12][5] ), .I1(\i11/fifo_inst/buff[14][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3816.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3817 (.I0(\i11/fifo_inst/buff[15][5] ), .I1(\i11/fifo_inst/buff[13][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3817.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3818 (.I0(n2359), .I1(n2358), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1853), .O(n2360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3818.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3819 (.I0(\i11/fifo_inst/buff[4][5] ), .I1(\i11/fifo_inst/buff[6][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3819.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3820 (.I0(\i11/fifo_inst/buff[7][5] ), .I1(\i11/fifo_inst/buff[5][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3820.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3821 (.I0(n2362), .I1(n2361), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n2363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3821.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3822 (.I0(\i11/fifo_inst/buff[8][5] ), .I1(\i11/fifo_inst/buff[10][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3822.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3823 (.I0(\i11/fifo_inst/buff[11][5] ), .I1(\i11/fifo_inst/buff[9][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3823.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3824 (.I0(n2365), .I1(n2364), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3824.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3825 (.I0(n2357), .I1(n2360), .I2(n2363), .I3(n2366), 
            .O(n2367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3825.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3826 (.I0(\i11/fifo_inst/buff[20][5] ), .I1(\i11/fifo_inst/buff[22][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3826.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3827 (.I0(\i11/fifo_inst/buff[23][5] ), .I1(\i11/fifo_inst/buff[21][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3827.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3828 (.I0(n2369), .I1(n2368), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n2370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3828.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3829 (.I0(\i11/fifo_inst/buff[28][5] ), .I1(\i11/fifo_inst/buff[30][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3829.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3830 (.I0(\i11/fifo_inst/buff[31][5] ), .I1(\i11/fifo_inst/buff[29][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3830.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3831 (.I0(n2372), .I1(n2371), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1853), .O(n2373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3831.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3832 (.I0(\i11/fifo_inst/buff[16][5] ), .I1(\i11/fifo_inst/buff[18][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3832.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3833 (.I0(\i11/fifo_inst/buff[19][5] ), .I1(\i11/fifo_inst/buff[17][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3833.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3834 (.I0(n2375), .I1(n2374), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3834.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3835 (.I0(\i11/fifo_inst/buff[24][5] ), .I1(\i11/fifo_inst/buff[26][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3835.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3836 (.I0(\i11/fifo_inst/buff[27][5] ), .I1(\i11/fifo_inst/buff[25][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3836.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3837 (.I0(n2378), .I1(n2377), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3837.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3838 (.I0(n2370), .I1(n2373), .I2(n2376), .I3(n2379), 
            .O(n2380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3838.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3839 (.I0(n2380), .I1(n2367), .I2(n1882), .I3(n2246), 
            .O(n2381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3839.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3840 (.I0(n1780), .I1(\rx_d[5] ), .I2(n2381), .O(n2382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__3840.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__3841 (.I0(n2331), .I1(n1895), .I2(n2354), .I3(n2382), 
            .O(\fifo_inst/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4ff */ ;
    defparam LUT__3841.LUTMASK = 16'hf4ff;
    EFX_LUT4 LUT__3842 (.I0(\i11/fifo_inst/buff[84][6] ), .I1(\i11/fifo_inst/buff[86][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3842.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3843 (.I0(\i11/fifo_inst/buff[87][6] ), .I1(\i11/fifo_inst/buff[85][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2383), .O(n2384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3843.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3844 (.I0(\i11/fifo_inst/buff[116][6] ), .I1(\i11/fifo_inst/buff[118][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3844.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3845 (.I0(\i11/fifo_inst/buff[119][6] ), .I1(\i11/fifo_inst/buff[117][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2385), .O(n2386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3845.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3846 (.I0(n2386), .I1(n2384), .I2(n1785), .I3(n1881), 
            .O(n2387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3846.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3847 (.I0(\i11/fifo_inst/buff[80][6] ), .I1(\i11/fifo_inst/buff[82][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3847.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3848 (.I0(\i11/fifo_inst/buff[83][6] ), .I1(\i11/fifo_inst/buff[81][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2388), .O(n2389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3848.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3849 (.I0(\i11/fifo_inst/buff[112][6] ), .I1(\i11/fifo_inst/buff[114][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3849.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3850 (.I0(\i11/fifo_inst/buff[115][6] ), .I1(\i11/fifo_inst/buff[113][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2390), .O(n2391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3850.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3851 (.I0(n2391), .I1(n2389), .I2(n1881), .I3(n1785), 
            .O(n2392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3851.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3852 (.I0(n2387), .I1(n2392), .I2(n1795), .O(n2393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3852.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3853 (.I0(\i11/fifo_inst/buff[92][6] ), .I1(\i11/fifo_inst/buff[94][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3853.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3854 (.I0(\i11/fifo_inst/buff[95][6] ), .I1(\i11/fifo_inst/buff[93][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2394), .O(n2395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3854.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3855 (.I0(\i11/fifo_inst/buff[124][6] ), .I1(\i11/fifo_inst/buff[126][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3855.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3856 (.I0(\i11/fifo_inst/buff[127][6] ), .I1(\i11/fifo_inst/buff[125][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2396), .O(n2397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3856.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3857 (.I0(n2397), .I1(n2395), .I2(n1785), .I3(n1881), 
            .O(n2398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3857.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3858 (.I0(\i11/fifo_inst/buff[88][6] ), .I1(\i11/fifo_inst/buff[90][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3858.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3859 (.I0(\i11/fifo_inst/buff[91][6] ), .I1(\i11/fifo_inst/buff[89][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2399), .O(n2400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3859.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3860 (.I0(\i11/fifo_inst/buff[120][6] ), .I1(\i11/fifo_inst/buff[122][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3860.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3861 (.I0(\i11/fifo_inst/buff[123][6] ), .I1(\i11/fifo_inst/buff[121][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2401), .O(n2402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3861.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3862 (.I0(n2402), .I1(n2400), .I2(n1881), .I3(n1785), 
            .O(n2403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3862.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3863 (.I0(n2398), .I1(n2403), .I2(n1795), .O(n2404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__3863.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__3864 (.I0(\i11/fifo_inst/buff[68][6] ), .I1(\i11/fifo_inst/buff[70][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3864.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3865 (.I0(\i11/fifo_inst/buff[71][6] ), .I1(\i11/fifo_inst/buff[69][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3865.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3866 (.I0(n2406), .I1(n2405), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n2407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3866.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3867 (.I0(\i11/fifo_inst/buff[76][6] ), .I1(\i11/fifo_inst/buff[78][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3867.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3868 (.I0(\i11/fifo_inst/buff[79][6] ), .I1(\i11/fifo_inst/buff[77][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3868.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3869 (.I0(n2409), .I1(n2408), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1853), .O(n2410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3869.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3870 (.I0(\i11/fifo_inst/buff[64][6] ), .I1(\i11/fifo_inst/buff[66][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3870.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3871 (.I0(\i11/fifo_inst/buff[67][6] ), .I1(\i11/fifo_inst/buff[65][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3871.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3872 (.I0(n2412), .I1(n2411), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3872.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3873 (.I0(\i11/fifo_inst/buff[72][6] ), .I1(\i11/fifo_inst/buff[74][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3873.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3874 (.I0(\i11/fifo_inst/buff[75][6] ), .I1(\i11/fifo_inst/buff[73][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3874.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3875 (.I0(n2415), .I1(n2414), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3875.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3876 (.I0(n2407), .I1(n2410), .I2(n2413), .I3(n2416), 
            .O(n2417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3876.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3877 (.I0(\i11/fifo_inst/buff[100][6] ), .I1(\i11/fifo_inst/buff[102][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3877.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3878 (.I0(\i11/fifo_inst/buff[103][6] ), .I1(\i11/fifo_inst/buff[101][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3878.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3879 (.I0(n2419), .I1(n2418), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n2420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3879.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3880 (.I0(\i11/fifo_inst/buff[108][6] ), .I1(\i11/fifo_inst/buff[110][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3880.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3881 (.I0(\i11/fifo_inst/buff[111][6] ), .I1(\i11/fifo_inst/buff[109][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3881.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3882 (.I0(n2422), .I1(n2421), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1853), .O(n2423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3882.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3883 (.I0(\i11/fifo_inst/buff[96][6] ), .I1(\i11/fifo_inst/buff[98][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3883.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3884 (.I0(\i11/fifo_inst/buff[99][6] ), .I1(\i11/fifo_inst/buff[97][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3884.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3885 (.I0(n2425), .I1(n2424), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3885.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3886 (.I0(\i11/fifo_inst/buff[104][6] ), .I1(\i11/fifo_inst/buff[106][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3886.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3887 (.I0(\i11/fifo_inst/buff[107][6] ), .I1(\i11/fifo_inst/buff[105][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3887.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3888 (.I0(n2428), .I1(n2427), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3888.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3889 (.I0(n2420), .I1(n2423), .I2(n2426), .I3(n2429), 
            .O(n2430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3889.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3890 (.I0(n2430), .I1(n2417), .I2(n1881), .O(n2431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3890.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3891 (.I0(n2404), .I1(n2393), .I2(n2431), .I3(n1882), 
            .O(n2432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3891.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3892 (.I0(n1780), .I1(\rx_d[6] ), .O(n2433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3892.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3893 (.I0(\i11/fifo_inst/buff[24][6] ), .I1(\i11/fifo_inst/buff[26][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3893.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3894 (.I0(\i11/fifo_inst/buff[27][6] ), .I1(\i11/fifo_inst/buff[25][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2434), .O(n2435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3894.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3895 (.I0(\i11/fifo_inst/buff[8][6] ), .I1(\i11/fifo_inst/buff[10][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3895.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3896 (.I0(\i11/fifo_inst/buff[11][6] ), .I1(\i11/fifo_inst/buff[9][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2436), .O(n2437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3896.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3897 (.I0(n2437), .I1(n2435), .I2(\fifo_inst/rd_index[4] ), 
            .I3(n1785), .O(n2438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__3897.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__3898 (.I0(\i11/fifo_inst/buff[12][6] ), .I1(\i11/fifo_inst/buff[14][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3898.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3899 (.I0(\i11/fifo_inst/buff[15][6] ), .I1(\i11/fifo_inst/buff[13][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2439), .O(n2440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3899.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3900 (.I0(\i11/fifo_inst/buff[28][6] ), .I1(\i11/fifo_inst/buff[30][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3900.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3901 (.I0(\i11/fifo_inst/buff[31][6] ), .I1(\i11/fifo_inst/buff[29][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2441), .O(n2442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3901.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3902 (.I0(n2442), .I1(n2440), .I2(n1785), .I3(\fifo_inst/rd_index[4] ), 
            .O(n2443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3902.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3903 (.I0(n1795), .I1(n2438), .I2(n2443), .I3(n1881), 
            .O(n2444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__3903.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__3904 (.I0(\i11/fifo_inst/buff[23][6] ), .I1(\i11/fifo_inst/buff[21][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3904.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3905 (.I0(\i11/fifo_inst/buff[20][6] ), .I1(\i11/fifo_inst/buff[22][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3905.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3906 (.I0(\i11/fifo_inst/buff[16][6] ), .I1(\i11/fifo_inst/buff[18][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3906.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3907 (.I0(\i11/fifo_inst/buff[19][6] ), .I1(\i11/fifo_inst/buff[17][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2447), .O(n2448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3907.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3908 (.I0(n2446), .I1(n2445), .I2(n2448), .I3(n1785), 
            .O(n2449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__3908.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__3909 (.I0(\i11/fifo_inst/buff[7][6] ), .I1(\i11/fifo_inst/buff[5][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3909.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3910 (.I0(\i11/fifo_inst/buff[4][6] ), .I1(\i11/fifo_inst/buff[6][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3910.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3911 (.I0(\i11/fifo_inst/buff[0][6] ), .I1(\i11/fifo_inst/buff[2][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3911.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3912 (.I0(\i11/fifo_inst/buff[3][6] ), .I1(\i11/fifo_inst/buff[1][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2452), .O(n2453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3912.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3913 (.I0(n2451), .I1(n2450), .I2(n2453), .I3(n1785), 
            .O(n2454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__3913.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__3914 (.I0(n2454), .I1(n2449), .I2(n1882), .I3(n1795), 
            .O(n2455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3914.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3915 (.I0(\i11/fifo_inst/buff[52][6] ), .I1(\i11/fifo_inst/buff[54][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3915.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3916 (.I0(\i11/fifo_inst/buff[55][6] ), .I1(\i11/fifo_inst/buff[53][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3916.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3917 (.I0(\i11/fifo_inst/buff[48][6] ), .I1(\i11/fifo_inst/buff[50][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3917.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3918 (.I0(\i11/fifo_inst/buff[51][6] ), .I1(\i11/fifo_inst/buff[49][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2458), .O(n2459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3918.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3919 (.I0(n2457), .I1(n2456), .I2(n2459), .I3(n1785), 
            .O(n2460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3919.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3920 (.I0(\i11/fifo_inst/buff[59][6] ), .I1(\i11/fifo_inst/buff[57][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3920.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__3921 (.I0(\i11/fifo_inst/buff[56][6] ), .I1(\i11/fifo_inst/buff[58][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3921.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3922 (.I0(\i11/fifo_inst/buff[60][6] ), .I1(\i11/fifo_inst/buff[62][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3922.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3923 (.I0(\i11/fifo_inst/buff[63][6] ), .I1(\i11/fifo_inst/buff[61][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2463), .O(n2464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3923.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3924 (.I0(n2462), .I1(n2461), .I2(n2464), .I3(n1785), 
            .O(n2465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__3924.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__3925 (.I0(n2465), .I1(n2460), .I2(n1795), .I3(n1829), 
            .O(n2466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__3925.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__3926 (.I0(\i11/fifo_inst/buff[44][6] ), .I1(\i11/fifo_inst/buff[46][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3926.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3927 (.I0(\i11/fifo_inst/buff[47][6] ), .I1(\i11/fifo_inst/buff[45][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2467), .O(n2468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3927.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3928 (.I0(\i11/fifo_inst/buff[40][6] ), .I1(\i11/fifo_inst/buff[42][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3928.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3929 (.I0(\i11/fifo_inst/buff[43][6] ), .I1(\i11/fifo_inst/buff[41][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3929.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3930 (.I0(n2470), .I1(n2469), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3930.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3931 (.I0(\i11/fifo_inst/buff[36][6] ), .I1(\i11/fifo_inst/buff[38][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3931.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3932 (.I0(\i11/fifo_inst/buff[39][6] ), .I1(\i11/fifo_inst/buff[37][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3932.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3933 (.I0(n2473), .I1(n2472), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n2474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3933.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3934 (.I0(\i11/fifo_inst/buff[32][6] ), .I1(\i11/fifo_inst/buff[34][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3934.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3935 (.I0(\i11/fifo_inst/buff[35][6] ), .I1(\i11/fifo_inst/buff[33][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3935.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3936 (.I0(n2476), .I1(n2475), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3936.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3937 (.I0(n1794), .I1(n2471), .I2(n2474), .I3(n2477), 
            .O(n2478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3937.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3938 (.I0(n2468), .I1(n1853), .I2(n2478), .I3(n1838), 
            .O(n2479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__3938.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__3939 (.I0(n2455), .I1(n2444), .I2(n2466), .I3(n2479), 
            .O(n2480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__3939.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__3940 (.I0(n2432), .I1(n1895), .I2(n2433), .I3(n2480), 
            .O(\fifo_inst/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__3940.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__3941 (.I0(\i11/fifo_inst/buff[84][7] ), .I1(\i11/fifo_inst/buff[86][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3941.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3942 (.I0(\i11/fifo_inst/buff[87][7] ), .I1(\i11/fifo_inst/buff[85][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2481), .O(n2482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3942.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3943 (.I0(\i11/fifo_inst/buff[116][7] ), .I1(\i11/fifo_inst/buff[118][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3943.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3944 (.I0(\i11/fifo_inst/buff[119][7] ), .I1(\i11/fifo_inst/buff[117][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2483), .O(n2484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3944.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3945 (.I0(n2484), .I1(n2482), .I2(n1785), .I3(n1881), 
            .O(n2485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3945.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3946 (.I0(\i11/fifo_inst/buff[80][7] ), .I1(\i11/fifo_inst/buff[82][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3946.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3947 (.I0(\i11/fifo_inst/buff[83][7] ), .I1(\i11/fifo_inst/buff[81][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2486), .O(n2487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3947.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3948 (.I0(\i11/fifo_inst/buff[112][7] ), .I1(\i11/fifo_inst/buff[114][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3948.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3949 (.I0(\i11/fifo_inst/buff[115][7] ), .I1(\i11/fifo_inst/buff[113][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2488), .O(n2489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3949.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3950 (.I0(n2489), .I1(n2487), .I2(n1881), .I3(n1785), 
            .O(n2490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3950.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3951 (.I0(n2485), .I1(n2490), .I2(n1795), .O(n2491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3951.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3952 (.I0(\i11/fifo_inst/buff[92][7] ), .I1(\i11/fifo_inst/buff[94][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3952.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3953 (.I0(\i11/fifo_inst/buff[95][7] ), .I1(\i11/fifo_inst/buff[93][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2492), .O(n2493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3953.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3954 (.I0(\i11/fifo_inst/buff[124][7] ), .I1(\i11/fifo_inst/buff[126][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3954.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3955 (.I0(\i11/fifo_inst/buff[127][7] ), .I1(\i11/fifo_inst/buff[125][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2494), .O(n2495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3955.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3956 (.I0(n2495), .I1(n2493), .I2(n1785), .I3(n1881), 
            .O(n2496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3956.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3957 (.I0(\i11/fifo_inst/buff[88][7] ), .I1(\i11/fifo_inst/buff[90][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3957.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3958 (.I0(\i11/fifo_inst/buff[91][7] ), .I1(\i11/fifo_inst/buff[89][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2497), .O(n2498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3958.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3959 (.I0(\i11/fifo_inst/buff[120][7] ), .I1(\i11/fifo_inst/buff[122][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__3959.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__3960 (.I0(\i11/fifo_inst/buff[123][7] ), .I1(\i11/fifo_inst/buff[121][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2499), .O(n2500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__3960.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__3961 (.I0(n2500), .I1(n2498), .I2(n1881), .I3(n1785), 
            .O(n2501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3961.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3962 (.I0(n2496), .I1(n2501), .I2(n1795), .O(n2502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__3962.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__3963 (.I0(\i11/fifo_inst/buff[76][7] ), .I1(\i11/fifo_inst/buff[78][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3963.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3964 (.I0(\i11/fifo_inst/buff[79][7] ), .I1(\i11/fifo_inst/buff[77][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3964.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3965 (.I0(n2504), .I1(n2503), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1853), .O(n2505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3965.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3966 (.I0(\i11/fifo_inst/buff[72][7] ), .I1(\i11/fifo_inst/buff[74][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3966.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3967 (.I0(\i11/fifo_inst/buff[75][7] ), .I1(\i11/fifo_inst/buff[73][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3967.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3968 (.I0(n2507), .I1(n2506), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3968.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3969 (.I0(\i11/fifo_inst/buff[68][7] ), .I1(\i11/fifo_inst/buff[70][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3969.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3970 (.I0(\i11/fifo_inst/buff[71][7] ), .I1(\i11/fifo_inst/buff[69][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3970.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3971 (.I0(n2510), .I1(n2509), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n2511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3971.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3972 (.I0(\i11/fifo_inst/buff[64][7] ), .I1(\i11/fifo_inst/buff[66][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3972.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3973 (.I0(\i11/fifo_inst/buff[67][7] ), .I1(\i11/fifo_inst/buff[65][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3973.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3974 (.I0(n2513), .I1(n2512), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3974.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3975 (.I0(n2505), .I1(n2508), .I2(n2511), .I3(n2514), 
            .O(n2515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3975.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3976 (.I0(\i11/fifo_inst/buff[96][7] ), .I1(\i11/fifo_inst/buff[98][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3976.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3977 (.I0(\i11/fifo_inst/buff[99][7] ), .I1(\i11/fifo_inst/buff[97][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3977.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3978 (.I0(n2517), .I1(n2516), .I2(n1857), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3978.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3979 (.I0(\i11/fifo_inst/buff[108][7] ), .I1(\i11/fifo_inst/buff[110][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3979.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3980 (.I0(\i11/fifo_inst/buff[111][7] ), .I1(\i11/fifo_inst/buff[109][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3980.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3981 (.I0(n2520), .I1(n2519), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1853), .O(n2521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3981.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3982 (.I0(\i11/fifo_inst/buff[100][7] ), .I1(\i11/fifo_inst/buff[102][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3982.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3983 (.I0(\i11/fifo_inst/buff[103][7] ), .I1(\i11/fifo_inst/buff[101][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3983.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3984 (.I0(n2523), .I1(n2522), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n2524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__3984.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__3985 (.I0(\i11/fifo_inst/buff[104][7] ), .I1(\i11/fifo_inst/buff[106][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3985.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3986 (.I0(\i11/fifo_inst/buff[107][7] ), .I1(\i11/fifo_inst/buff[105][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3986.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3987 (.I0(n2526), .I1(n2525), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__3987.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__3988 (.I0(n2518), .I1(n2521), .I2(n2524), .I3(n2527), 
            .O(n2528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3988.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3989 (.I0(n2528), .I1(n2515), .I2(n1881), .O(n2529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3989.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3990 (.I0(n2502), .I1(n2491), .I2(n2529), .I3(n1882), 
            .O(n2530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3990.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3991 (.I0(n1780), .I1(\rx_d[7] ), .O(n2531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3991.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3992 (.I0(\i11/fifo_inst/buff[12][7] ), .I1(\i11/fifo_inst/buff[14][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__3992.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__3993 (.I0(\i11/fifo_inst/buff[15][7] ), .I1(\i11/fifo_inst/buff[13][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2532), .O(n2533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__3993.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__3994 (.I0(\i11/fifo_inst/buff[28][7] ), .I1(\i11/fifo_inst/buff[30][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__3994.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__3995 (.I0(\i11/fifo_inst/buff[31][7] ), .I1(\i11/fifo_inst/buff[29][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__3995.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__3996 (.I0(n2535), .I1(n2534), .I2(\fifo_inst/rd_index[4] ), 
            .I3(n1785), .O(n2536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__3996.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__3997 (.I0(\fifo_inst/rd_index[4] ), .I1(n2533), .I2(n2532), 
            .I3(n2536), .O(n2537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbe00 */ ;
    defparam LUT__3997.LUTMASK = 16'hbe00;
    EFX_LUT4 LUT__3998 (.I0(\i11/fifo_inst/buff[8][7] ), .I1(\i11/fifo_inst/buff[10][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__3998.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__3999 (.I0(\i11/fifo_inst/buff[11][7] ), .I1(\i11/fifo_inst/buff[9][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__3999.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4000 (.I0(\i11/fifo_inst/buff[27][7] ), .I1(\i11/fifo_inst/buff[25][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4000.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4001 (.I0(\i11/fifo_inst/buff[24][7] ), .I1(\i11/fifo_inst/buff[26][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4001.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4002 (.I0(n2541), .I1(n2540), .I2(\fifo_inst/rd_index[4] ), 
            .I3(n1785), .O(n2542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__4002.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__4003 (.I0(n2538), .I1(n2539), .I2(\fifo_inst/rd_index[4] ), 
            .I3(n2542), .O(n2543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__4003.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__4004 (.I0(n1795), .I1(n2537), .I2(n2543), .I3(n1881), 
            .O(n2544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__4004.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__4005 (.I0(\i11/fifo_inst/buff[7][7] ), .I1(\i11/fifo_inst/buff[5][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4005.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4006 (.I0(\i11/fifo_inst/buff[4][7] ), .I1(\i11/fifo_inst/buff[6][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4006.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4007 (.I0(\i11/fifo_inst/buff[20][7] ), .I1(\i11/fifo_inst/buff[22][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__4007.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__4008 (.I0(\i11/fifo_inst/buff[23][7] ), .I1(\i11/fifo_inst/buff[21][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2547), .O(n2548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__4008.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__4009 (.I0(n2546), .I1(n2545), .I2(n2548), .I3(n1882), 
            .O(n2549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__4009.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__4010 (.I0(\i11/fifo_inst/buff[0][7] ), .I1(\i11/fifo_inst/buff[2][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__4010.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__4011 (.I0(\i11/fifo_inst/buff[3][7] ), .I1(\i11/fifo_inst/buff[1][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2550), .O(n2551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__4011.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__4012 (.I0(\i11/fifo_inst/buff[16][7] ), .I1(\i11/fifo_inst/buff[18][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__4012.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__4013 (.I0(\i11/fifo_inst/buff[19][7] ), .I1(\i11/fifo_inst/buff[17][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2552), .O(n2553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__4013.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__4014 (.I0(n2553), .I1(n2551), .I2(n1882), .I3(n1785), 
            .O(n2554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__4014.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__4015 (.I0(n2549), .I1(n1785), .I2(n2554), .I3(n1795), 
            .O(n2555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__4015.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__4016 (.I0(\i11/fifo_inst/buff[52][7] ), .I1(\i11/fifo_inst/buff[54][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4016.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4017 (.I0(\i11/fifo_inst/buff[55][7] ), .I1(\i11/fifo_inst/buff[53][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4017.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4018 (.I0(\i11/fifo_inst/buff[48][7] ), .I1(\i11/fifo_inst/buff[50][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4018.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4019 (.I0(\i11/fifo_inst/buff[51][7] ), .I1(\i11/fifo_inst/buff[49][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2558), .O(n2559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4019.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4020 (.I0(n2557), .I1(n2556), .I2(n2559), .I3(n1785), 
            .O(n2560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__4020.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__4021 (.I0(\i11/fifo_inst/buff[59][7] ), .I1(\i11/fifo_inst/buff[57][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__4021.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__4022 (.I0(\i11/fifo_inst/buff[56][7] ), .I1(\i11/fifo_inst/buff[58][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__4022.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__4023 (.I0(\i11/fifo_inst/buff[60][7] ), .I1(\i11/fifo_inst/buff[62][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4023.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4024 (.I0(\i11/fifo_inst/buff[63][7] ), .I1(\i11/fifo_inst/buff[61][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2563), .O(n2564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4024.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4025 (.I0(n2562), .I1(n2561), .I2(n2564), .I3(n1785), 
            .O(n2565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__4025.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__4026 (.I0(n2565), .I1(n2560), .I2(n1795), .I3(n1829), 
            .O(n2566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__4026.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__4027 (.I0(\i11/fifo_inst/buff[36][7] ), .I1(\i11/fifo_inst/buff[38][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4027.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4028 (.I0(\i11/fifo_inst/buff[39][7] ), .I1(\i11/fifo_inst/buff[37][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4028.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4029 (.I0(n2568), .I1(n2567), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n1861), .O(n2569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__4029.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__4030 (.I0(\i11/fifo_inst/buff[32][7] ), .I1(\i11/fifo_inst/buff[34][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__4030.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__4031 (.I0(\i11/fifo_inst/buff[35][7] ), .I1(\i11/fifo_inst/buff[33][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n2570), .O(n2571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__4031.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__4032 (.I0(n1857), .I1(n2571), .I2(n1794), .O(n2572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__4032.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__4033 (.I0(\i11/fifo_inst/buff[47][7] ), .I1(\i11/fifo_inst/buff[45][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n2573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__4033.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__4034 (.I0(\i11/fifo_inst/buff[44][7] ), .I1(\i11/fifo_inst/buff[46][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__4034.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__4035 (.I0(\i11/fifo_inst/buff[40][7] ), .I1(\i11/fifo_inst/buff[42][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4035.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4036 (.I0(\i11/fifo_inst/buff[43][7] ), .I1(\i11/fifo_inst/buff[41][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n2576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__4036.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__4037 (.I0(n2576), .I1(n2575), .I2(n1865), .I3(\fifo_inst/rd_index[0] ), 
            .O(n2577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__4037.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__4038 (.I0(n2574), .I1(n2573), .I2(n1853), .I3(n2577), 
            .O(n2578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__4038.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__4039 (.I0(n2569), .I1(n2578), .I2(n2572), .I3(n1838), 
            .O(n2579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__4039.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__4040 (.I0(n2555), .I1(n2544), .I2(n2566), .I3(n2579), 
            .O(n2580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__4040.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__4041 (.I0(n2530), .I1(n1895), .I2(n2531), .I3(n2580), 
            .O(\fifo_inst/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__4041.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__4042 (.I0(n1751), .I1(n1748), .O(\i11/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4042.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4043 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[2] ), 
            .O(n2581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4043.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4044 (.I0(\fifo_inst/wr_index[3] ), .I1(\fifo_inst/wr_index[4] ), 
            .I2(n1747), .I3(n2581), .O(\i11/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__4044.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__4045 (.I0(\fifo_inst/wr_index[3] ), .I1(\fifo_inst/wr_index[4] ), 
            .I2(n1751), .I3(n2581), .O(\i11/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__4045.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__4046 (.I0(\fifo_inst/wr_index[4] ), .I1(\fifo_inst/wr_index[3] ), 
            .O(n2582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__4046.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__4047 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[2] ), 
            .I2(n2582), .O(n2583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4047.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4048 (.I0(n1747), .I1(n2583), .O(\i11/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4048.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4049 (.I0(n1751), .I1(n2583), .O(\i11/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4049.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4050 (.I0(\fifo_inst/wr_index[2] ), .I1(\fifo_inst/wr_index[1] ), 
            .I2(n2582), .O(n2584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4050.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4051 (.I0(n1747), .I1(n2584), .O(\i11/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4051.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4052 (.I0(n1751), .I1(n2584), .O(\i11/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4052.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4053 (.I0(\fifo_inst/wr_index[1] ), .I1(n2582), .I2(\fifo_inst/wr_index[2] ), 
            .O(n2585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4053.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4054 (.I0(n1747), .I1(n2585), .O(\i11/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4054.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4055 (.I0(n1751), .I1(n2585), .O(\i11/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4055.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4056 (.I0(n1747), .I1(n2581), .I2(n2582), .O(\i11/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4056.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4057 (.I0(n1751), .I1(n2581), .I2(n2582), .O(\i11/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4057.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4058 (.I0(\fifo_inst/wr_index[3] ), .I1(\fifo_inst/wr_index[4] ), 
            .O(n2586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__4058.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__4059 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[2] ), 
            .I2(n2586), .O(n2587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4059.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4060 (.I0(n1747), .I1(n2587), .O(\i11/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4060.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4061 (.I0(n1751), .I1(n2587), .O(\i11/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4061.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4062 (.I0(\fifo_inst/wr_index[2] ), .I1(\fifo_inst/wr_index[1] ), 
            .I2(n2586), .O(n2588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4062.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4063 (.I0(n1747), .I1(n2588), .O(\i11/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4063.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4064 (.I0(n1751), .I1(n2588), .O(\i11/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4064.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4065 (.I0(\fifo_inst/wr_index[1] ), .I1(n2586), .I2(\fifo_inst/wr_index[2] ), 
            .O(n2589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4065.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4066 (.I0(n1747), .I1(n2589), .O(\i11/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4066.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4067 (.I0(n1751), .I1(n2589), .O(\i11/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4067.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4068 (.I0(n1747), .I1(n2581), .I2(n2586), .O(\i11/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4068.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4069 (.I0(n1751), .I1(n2581), .I2(n2586), .O(\i11/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4069.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4070 (.I0(\fifo_inst/wr_index[3] ), .I1(\fifo_inst/wr_index[4] ), 
            .O(n2590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4070.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4071 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[2] ), 
            .I2(n2590), .O(n2591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4071.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4072 (.I0(n1747), .I1(n2591), .O(\i11/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4072.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4073 (.I0(n1751), .I1(n2591), .O(\i11/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4073.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4074 (.I0(\fifo_inst/wr_index[2] ), .I1(\fifo_inst/wr_index[1] ), 
            .I2(n2590), .O(n2592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4074.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4075 (.I0(n1747), .I1(n2592), .O(\i11/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4075.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4076 (.I0(n1751), .I1(n2592), .O(\i11/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4076.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4077 (.I0(\fifo_inst/wr_index[1] ), .I1(n2590), .I2(\fifo_inst/wr_index[2] ), 
            .O(n2593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4077.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4078 (.I0(n1747), .I1(n2593), .O(\i11/n104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4078.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4079 (.I0(n1751), .I1(n2593), .O(\i11/n103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4079.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4080 (.I0(n1747), .I1(n2581), .I2(n2590), .O(\i11/n102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4080.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4081 (.I0(n1751), .I1(n2581), .I2(n2590), .O(\i11/n101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4081.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4082 (.I0(\fifo_inst/wr_index[6] ), .I1(\fifo_inst/wr_index[5] ), 
            .I2(n1746), .O(n2594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4082.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4083 (.I0(n2594), .I1(n1752), .O(\i11/n100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4083.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4084 (.I0(\fifo_inst/wr_index[6] ), .I1(\fifo_inst/wr_index[5] ), 
            .I2(n1750), .O(n2595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4084.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4085 (.I0(n2595), .I1(n1752), .O(\i11/n99 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4085.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4086 (.I0(n2594), .I1(n1749), .O(\i11/n98 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4086.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4087 (.I0(n2595), .I1(n1749), .O(\i11/n97 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4087.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4088 (.I0(n2594), .I1(n1748), .O(\i11/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4088.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4089 (.I0(n2595), .I1(n1748), .O(\i11/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4089.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4090 (.I0(\fifo_inst/wr_index[0] ), .I1(\fifo_inst/wr_index[7] ), 
            .I2(n2581), .O(n2596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__4090.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__4091 (.I0(\fifo_inst/wr_index[6] ), .I1(\fifo_inst/wr_index[5] ), 
            .I2(n2596), .O(n2597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4091.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4092 (.I0(\fifo_inst/wr_index[3] ), .I1(\fifo_inst/wr_index[4] ), 
            .I2(n2597), .I3(n1745), .O(\i11/n94 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__4092.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__4093 (.I0(\fifo_inst/wr_index[7] ), .I1(\fifo_inst/wr_index[0] ), 
            .I2(n2581), .O(n2598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4093.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4094 (.I0(\fifo_inst/wr_index[6] ), .I1(\fifo_inst/wr_index[5] ), 
            .I2(n2598), .O(n2599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4094.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4095 (.I0(\fifo_inst/wr_index[3] ), .I1(\fifo_inst/wr_index[4] ), 
            .I2(n2599), .I3(n1745), .O(\i11/n93 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__4095.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__4096 (.I0(n2594), .I1(n2583), .O(\i11/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4096.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4097 (.I0(n2595), .I1(n2583), .O(\i11/n91 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4097.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4098 (.I0(n2594), .I1(n2584), .O(\i11/n90 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4098.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4099 (.I0(n2595), .I1(n2584), .O(\i11/n89 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4099.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4100 (.I0(n2594), .I1(n2585), .O(\i11/n88 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4100.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4101 (.I0(n2595), .I1(n2585), .O(\i11/n87 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4101.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4102 (.I0(n2597), .I1(n1745), .I2(n2582), .O(\i11/n86 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4102.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4103 (.I0(n2599), .I1(n1745), .I2(n2582), .O(\i11/n85 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4103.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4104 (.I0(n2594), .I1(n2587), .O(\i11/n84 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4104.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4105 (.I0(n2595), .I1(n2587), .O(\i11/n83 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4105.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4106 (.I0(n2594), .I1(n2588), .O(\i11/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4106.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4107 (.I0(n2595), .I1(n2588), .O(\i11/n81 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4107.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4108 (.I0(n2594), .I1(n2589), .O(\i11/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4108.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4109 (.I0(n2595), .I1(n2589), .O(\i11/n79 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4109.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4110 (.I0(n2597), .I1(n1745), .I2(n2586), .O(\i11/n78 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4110.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4111 (.I0(n2599), .I1(n1745), .I2(n2586), .O(\i11/n77 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4111.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4112 (.I0(n2594), .I1(n2591), .O(\i11/n76 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4112.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4113 (.I0(n2595), .I1(n2591), .O(\i11/n75 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4113.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4114 (.I0(n2594), .I1(n2592), .O(\i11/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4114.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4115 (.I0(n2595), .I1(n2592), .O(\i11/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4115.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4116 (.I0(n2594), .I1(n2593), .O(\i11/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4116.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4117 (.I0(n2595), .I1(n2593), .O(\i11/n71 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4117.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4118 (.I0(n2597), .I1(n1745), .I2(n2590), .O(\i11/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4118.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4119 (.I0(n2599), .I1(n1745), .I2(n2590), .O(\i11/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4119.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4120 (.I0(\fifo_inst/wr_index[5] ), .I1(n1746), .I2(\fifo_inst/wr_index[6] ), 
            .O(n2600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4120.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4121 (.I0(n2600), .I1(n1752), .O(\i11/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4121.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4122 (.I0(\fifo_inst/wr_index[5] ), .I1(n1750), .I2(\fifo_inst/wr_index[6] ), 
            .O(n2601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4122.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4123 (.I0(n2601), .I1(n1752), .O(\i11/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4123.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4124 (.I0(n2600), .I1(n1749), .O(\i11/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4124.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4125 (.I0(n2601), .I1(n1749), .O(\i11/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4125.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4126 (.I0(n2600), .I1(n1748), .O(\i11/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4126.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4127 (.I0(n2601), .I1(n1748), .O(\i11/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4127.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4128 (.I0(\fifo_inst/wr_index[5] ), .I1(n2596), .I2(\fifo_inst/wr_index[6] ), 
            .O(n2602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4128.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4129 (.I0(\fifo_inst/wr_index[3] ), .I1(\fifo_inst/wr_index[4] ), 
            .I2(n2602), .I3(n1745), .O(\i11/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__4129.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__4130 (.I0(\fifo_inst/wr_index[5] ), .I1(n2598), .I2(\fifo_inst/wr_index[6] ), 
            .O(n2603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__4130.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__4131 (.I0(\fifo_inst/wr_index[3] ), .I1(\fifo_inst/wr_index[4] ), 
            .I2(n2603), .I3(n1745), .O(\i11/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__4131.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__4132 (.I0(n2600), .I1(n2583), .O(\i11/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4132.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4133 (.I0(n2601), .I1(n2583), .O(\i11/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4133.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4134 (.I0(n2600), .I1(n2584), .O(\i11/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4134.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4135 (.I0(n2601), .I1(n2584), .O(\i11/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4135.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4136 (.I0(n2600), .I1(n2585), .O(\i11/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4136.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4137 (.I0(n2601), .I1(n2585), .O(\i11/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4137.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4138 (.I0(n2602), .I1(n1745), .I2(n2582), .O(\i11/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4138.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4139 (.I0(n2603), .I1(n1745), .I2(n2582), .O(\i11/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4139.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4140 (.I0(n2600), .I1(n2587), .O(\i11/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4140.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4141 (.I0(n2601), .I1(n2587), .O(\i11/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4141.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4142 (.I0(n2600), .I1(n2588), .O(\i11/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4142.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4143 (.I0(n2601), .I1(n2588), .O(\i11/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4143.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4144 (.I0(n2600), .I1(n2589), .O(\i11/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4144.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4145 (.I0(n2601), .I1(n2589), .O(\i11/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4145.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4146 (.I0(n2602), .I1(n1745), .I2(n2586), .O(\i11/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4146.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4147 (.I0(n2603), .I1(n1745), .I2(n2586), .O(\i11/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4147.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4148 (.I0(n2600), .I1(n2591), .O(\i11/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4148.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4149 (.I0(n2601), .I1(n2591), .O(\i11/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4149.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4150 (.I0(n2600), .I1(n2592), .O(\i11/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4150.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4151 (.I0(n2601), .I1(n2592), .O(\i11/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4151.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4152 (.I0(n2600), .I1(n2593), .O(\i11/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4152.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4153 (.I0(n2601), .I1(n2593), .O(\i11/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4153.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4154 (.I0(n2602), .I1(n1745), .I2(n2590), .O(\i11/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4154.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4155 (.I0(n2603), .I1(n1745), .I2(n2590), .O(\i11/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4155.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4156 (.I0(n1746), .I1(\fifo_inst/wr_index[5] ), .I2(\fifo_inst/wr_index[6] ), 
            .O(n2604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4156.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4157 (.I0(n2604), .I1(n1752), .O(\i11/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4157.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4158 (.I0(n1750), .I1(\fifo_inst/wr_index[5] ), .I2(\fifo_inst/wr_index[6] ), 
            .O(n2605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4158.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4159 (.I0(n2605), .I1(n1752), .O(\i11/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4159.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4160 (.I0(n2604), .I1(n1749), .O(\i11/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4160.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4161 (.I0(n2605), .I1(n1749), .O(\i11/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4161.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4162 (.I0(n2604), .I1(n1748), .O(\i11/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4162.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4163 (.I0(n2605), .I1(n1748), .O(\i11/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4163.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4164 (.I0(n2596), .I1(\fifo_inst/wr_index[5] ), .I2(\fifo_inst/wr_index[6] ), 
            .O(n2606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4164.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4165 (.I0(\fifo_inst/wr_index[3] ), .I1(\fifo_inst/wr_index[4] ), 
            .I2(n2606), .I3(n1745), .O(\i11/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__4165.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__4166 (.I0(n2598), .I1(\fifo_inst/wr_index[5] ), .I2(\fifo_inst/wr_index[6] ), 
            .O(n2607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4166.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4167 (.I0(\fifo_inst/wr_index[3] ), .I1(\fifo_inst/wr_index[4] ), 
            .I2(n2607), .I3(n1745), .O(\i11/n29 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__4167.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__4168 (.I0(n2604), .I1(n2583), .O(\i11/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4168.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4169 (.I0(n2605), .I1(n2583), .O(\i11/n27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4169.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4170 (.I0(n2604), .I1(n2584), .O(\i11/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4170.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4171 (.I0(n2605), .I1(n2584), .O(\i11/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4171.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4172 (.I0(n2604), .I1(n2585), .O(\i11/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4172.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4173 (.I0(n2605), .I1(n2585), .O(\i11/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4173.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4174 (.I0(n2606), .I1(n1745), .I2(n2582), .O(\i11/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4174.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4175 (.I0(n2607), .I1(n1745), .I2(n2582), .O(\i11/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4175.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4176 (.I0(n2604), .I1(n2587), .O(\i11/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4176.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4177 (.I0(n2605), .I1(n2587), .O(\i11/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4177.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4178 (.I0(n2604), .I1(n2588), .O(\i11/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4178.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4179 (.I0(n2605), .I1(n2588), .O(\i11/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4179.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4180 (.I0(n2604), .I1(n2589), .O(\i11/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4180.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4181 (.I0(n2605), .I1(n2589), .O(\i11/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4181.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4182 (.I0(n2606), .I1(n1745), .I2(n2586), .O(\i11/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4182.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4183 (.I0(n2607), .I1(n1745), .I2(n2586), .O(\i11/n13 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4183.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4184 (.I0(n2604), .I1(n2591), .O(\i11/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4184.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4185 (.I0(n2605), .I1(n2591), .O(\i11/n11 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4185.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4186 (.I0(n2604), .I1(n2592), .O(\i11/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4186.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4187 (.I0(n2605), .I1(n2592), .O(\i11/n9 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4187.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4188 (.I0(n2604), .I1(n2593), .O(\i11/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4188.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4189 (.I0(n2605), .I1(n2593), .O(\i11/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4189.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4190 (.I0(n2606), .I1(n1745), .I2(n2590), .O(\i11/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4190.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4191 (.I0(n2607), .I1(n1745), .I2(n2590), .O(\i11/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4191.LUTMASK = 16'h8080;
    EFX_LUT4 \tx_dac_fsm_inst/dctr[4]~FF_frt_0_rtinv  (.I0(\tx_dac_fsm_inst/dctr[4]~FF_frt_0_q_pinv ), 
            .O(\tx_dac_fsm_inst/dctr[4]~FF_frt_0_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \tx_dac_fsm_inst/dctr[4]~FF_frt_0_rtinv .LUTMASK = 16'h5555;
    EFX_GBUFCE CLKBUF__1 (.CE(1'b1), .I(tx_slowclk), .O(\tx_slowclk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__1.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(pll_clk), .O(\pll_clk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__tx_dac_fsm_inst/add_18/i2  (.I0(\tx_dac_fsm_inst/sym_ctr[0] ), 
            .I1(1'b1), .CI(1'b0), .CO(n2612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(95)
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/add_18/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/add_18/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__tx_dac_fsm_inst/sub_20/add_2/i4  (.I0(\tx_dac_fsm_inst/sym_ctr[2] ), 
            .I1(1'b1), .CI(1'b0), .CO(n2611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(97)
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/sub_20/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/sub_20/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__tx_dac_fsm_inst/sub_20/add_2/i5  (.I0(n1633), .I1(1'b1), 
            .CI(1'b0), .CO(n2610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(97)
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/sub_20/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/sub_20/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__tx_dac_fsm_inst/add_129/i4  (.I0(n1628), .I1(1'b1), 
            .CI(1'b0), .CO(n2609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(197)
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/add_129/i4 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/add_129/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__tx_dac_fsm_inst/add_136/i4  (.I0(n1617), .I1(1'b1), 
            .CI(1'b0), .CO(n2608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(208)
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/add_136/i4 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/add_136/i4 .I1_POLARITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dctr[1]~FF_frt_1  (.D(n1756), .CE(1'b1), .CLK(\tx_slowclk~O ), 
           .SR(reset_n), .Q(\tx_dac_fsm_inst/dctr[1]~FF_frt_1_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, INIT_VALUE=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(211)
    defparam \tx_dac_fsm_inst/dctr[1]~FF_frt_1 .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[1]~FF_frt_1 .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[1]~FF_frt_1 .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[1]~FF_frt_1 .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[1]~FF_frt_1 .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[1]~FF_frt_1 .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[1]~FF_frt_1 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dctr[4]~FF_frt_0  (.D(n1757), .CE(1'b1), .CLK(\tx_slowclk~O ), 
           .SR(reset_n), .Q(\tx_dac_fsm_inst/dctr[4]~FF_frt_0_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(211)
    defparam \tx_dac_fsm_inst/dctr[4]~FF_frt_0 .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[4]~FF_frt_0 .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[4]~FF_frt_0 .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[4]~FF_frt_0 .D_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[4]~FF_frt_0 .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[4]~FF_frt_0 .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[4]~FF_frt_0 .SR_SYNC_PRIORITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_beaf11be_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_beaf11be_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_beaf11be_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_beaf11be_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_beaf11be_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_beaf11be_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_beaf11be_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_beaf11be_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_beaf11be_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_beaf11be_0
// module not written out since it is a black box. 
//



//
// Verific Verilog Description of module WES207_top
//

module WES207_top (pll_clk, reset_n, tx_slowclk, led0, led1, SCLK, 
            SSB, MOSI, MISO, gpo_pins, lvds_tx_inst1_DATA);
    input pll_clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input reset_n /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input tx_slowclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output led0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output led1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input SCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input SSB /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MOSI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output MISO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]gpo_pins /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]lvds_tx_inst1_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    
    wire \reg_addr[4] , \reg_addr[3] , \spi_slave_inst/bitcnt[2] , \spi_slave_inst/bitcnt[1] , 
        \spi_slave_inst/sync_tx_en[1] , \reg_addr[2] , \reg_addr[1] , 
        \spi_slave_inst/bitcnt[0] , \spi_slave_inst/sync_mosi[1] , n19, 
        n20, rw_out, \reg_addr[0] , \spi_slave_inst/d_o[0] , \rx_d[0] , 
        addr_dv, rxdv, \spi_slave_inst/sync_sclk[0] , \spi_slave_inst/bitcnt[4] , 
        \reg_addr[5] , \spi_slave_inst/bitcnt[3] , \spi_slave_inst/sync_ss[0] , 
        \reg_addr[6] , \spi_slave_inst/d_o[1] , \spi_slave_inst/d_o[2] , 
        \spi_slave_inst/d_o[3] , \spi_slave_inst/d_o[4] , \spi_slave_inst/d_o[5] , 
        \spi_slave_inst/d_o[6] , \spi_slave_inst/d_o[7] , \rx_d[1] , \rx_d[2] , 
        \rx_d[3] , \rx_d[4] , \rx_d[5] , \rx_d[6] , \rx_d[7] , \spi_slave_inst/sync_sclk[1] , 
        \spi_slave_inst/sync_sclk[2] , \spi_slave_inst/sync_ss[1] , \spi_slave_inst/sync_ss[2] , 
        \data_from_led[7] , \data_from_led[6] , \data_from_led[5] , \data_from_led[4] , 
        \data_from_led[3] , \data_from_led[0] , \data_from_led[2] , \data_from_led[1] , 
        \led_inst/counter[0] , \led_inst/ctr_cfg_reg[0] , \led_inst/counter[1] , 
        \led_inst/counter[2] , \led_inst/counter[3] , \led_inst/counter[4] , 
        \led_inst/counter[5] , \led_inst/counter[6] , \led_inst/counter[7] , 
        \led_inst/counter[8] , \led_inst/counter[9] , \led_inst/counter[10] , 
        \led_inst/counter[11] , \led_inst/counter[12] , \led_inst/counter[13] , 
        \led_inst/counter[14] , \led_inst/counter[15] , \led_inst/counter[16] , 
        \led_inst/counter[17] , \led_inst/counter[18] , \led_inst/counter[19] , 
        \led_inst/counter[20] , \led_inst/counter[21] , \led_inst/counter[22] , 
        \led_inst/counter[23] , \led_inst/ctr_cfg_reg[1] , \led_inst/ctr_cfg_reg[2] , 
        \led_inst/ctr_cfg_reg[3] , \led_inst/ctr_cfg_reg[4] , \led_inst/ctr_cfg_reg[5] , 
        \led_inst/ctr_cfg_reg[6] , \led_inst/ctr_cfg_reg[7] , \gpo_inst/gp_config_reg[0] , 
        \gpo_inst/gp_config_reg[1] , \gpo_inst/gp_config_reg[2] , \gpo_inst/gp_config_reg[3] , 
        \gpo_inst/gp_config_reg[4] , \gpo_inst/gp_config_reg[5] , \gpo_inst/gp_config_reg[6] , 
        \gpo_inst/gp_config_reg[7] , \i14/fifo_inst/buff[3][2] , \i14/fifo_inst/buff[3][1] , 
        \i14/fifo_inst/buff[3][0] , \i14/fifo_inst/buff[2][7] , \tx_dac_fsm_inst/sym_ctr[0] , 
        \tx_dac_fsm_inst/sym_pos[0] , \tx_dac_fsm_inst/state_reg[0] , n109, 
        \tx_dac_fsm_inst/sym_ctr[1] , \tx_dac_fsm_inst/sym_ctr[2] , \tx_dac_fsm_inst/sym_ctr[3] , 
        n113, \i14/fifo_inst/buff[2][6] , n115, n116, \tx_dac_fsm_inst/zctr[0] , 
        n118, n119, \tx_dac_fsm_inst/sym_ctr[4] , n121, n122, \tx_dac_fsm_inst/dctr[0] , 
        n124, n125, \tx_dac_fsm_inst/dac_config_reg[0] , \tx_dac_fsm_inst/sym_pos[1] , 
        \tx_dac_fsm_inst/sym_pos[2] , \tx_dac_fsm_inst/sym_pos[3] , \tx_dac_fsm_inst/state_reg[1] , 
        \tx_dac_fsm_inst/state_reg[2] , \tx_dac_fsm_inst/state_reg[3] , 
        n133, n134, n135, n136, \tx_dac_fsm_inst/zctr[1] , \tx_dac_fsm_inst/zctr[2] , 
        \tx_dac_fsm_inst/zctr[3] , \tx_dac_fsm_inst/zctr[4] , \tx_dac_fsm_inst/zctr[5] , 
        \tx_dac_fsm_inst/dctr[1] , \tx_dac_fsm_inst/dctr[2] , \tx_dac_fsm_inst/dctr[3] , 
        \tx_dac_fsm_inst/dctr[4] , \tx_dac_fsm_inst/dctr[5] , n147, n148, 
        \fifo_inst/wr_index[0] , \fifo_inst/rd_index[0] , \fifo_inst/length[0] , 
        \fifo_inst/sync_wr[0] , \fifo_inst/sync_rd[0] , \fifo_inst/buff_head[0] , 
        \fifo_inst/wr_index[1] , \fifo_inst/wr_index[2] , \fifo_inst/wr_index[3] , 
        \fifo_inst/wr_index[4] , \fifo_inst/wr_index[5] , \fifo_inst/wr_index[6] , 
        \fifo_inst/wr_index[7] , \fifo_inst/rd_index[1] , \fifo_inst/rd_index[2] , 
        \fifo_inst/rd_index[3] , \fifo_inst/rd_index[4] , \fifo_inst/rd_index[5] , 
        \fifo_inst/rd_index[6] , \fifo_inst/rd_index[7] , \fifo_inst/length[1] , 
        \fifo_inst/length[2] , \fifo_inst/length[3] , \fifo_inst/length[4] , 
        \fifo_inst/length[5] , \fifo_inst/length[6] , \fifo_inst/length[7] , 
        \fifo_inst/sync_wr[1] , \fifo_inst/sync_rd[1] , \i14/fifo_inst/buff[0][1] , 
        \i14/fifo_inst/buff[0][4] , \i14/fifo_inst/buff[0][7] , \i14/fifo_inst/buff[1][2] , 
        \i14/fifo_inst/buff[1][5] , \i14/fifo_inst/buff[2][0] , \i14/fifo_inst/buff[2][3] , 
        \i14/fifo_inst/buff[2][5] , \fifo_inst/buff_head[1] , \fifo_inst/buff_head[2] , 
        \fifo_inst/buff_head[3] , \fifo_inst/buff_head[4] , \fifo_inst/buff_head[5] , 
        \fifo_inst/buff_head[6] , \fifo_inst/buff_head[7] , n193, n194, 
        \tx_fifo/wr_index[0] , \tx_fifo/rd_index[0] , \tx_fifo/length[0] , 
        \tx_fifo/sync_wr[0] , \tx_fifo/sync_rd[0] , \tx_fifo/buff_head[0] , 
        \tx_fifo/wr_index[1] , \tx_fifo/wr_index[2] , \tx_fifo/wr_index[3] , 
        \tx_fifo/wr_index[4] , \tx_fifo/wr_index[5] , \tx_fifo/wr_index[6] , 
        \tx_fifo/wr_index[7] , \tx_fifo/rd_index[1] , \tx_fifo/rd_index[2] , 
        \tx_fifo/rd_index[3] , \tx_fifo/rd_index[4] , \tx_fifo/rd_index[5] , 
        \tx_fifo/rd_index[6] , \tx_fifo/rd_index[7] , \tx_fifo/length[1] , 
        \tx_fifo/length[2] , \tx_fifo/length[3] , \tx_fifo/length[4] , 
        \tx_fifo/length[5] , \tx_fifo/length[6] , \tx_fifo/length[7] , 
        \tx_fifo/sync_wr[1] , \tx_fifo/sync_rd[1] , \i14/fifo_inst/buff[0][0] , 
        \i14/fifo_inst/buff[0][3] , \i14/fifo_inst/buff[0][6] , \i14/fifo_inst/buff[1][1] , 
        \i14/fifo_inst/buff[1][4] , \i14/fifo_inst/buff[1][7] , \i14/fifo_inst/buff[2][2] , 
        \tx_fifo/buff_head[1] , \tx_fifo/buff_head[2] , \tx_fifo/buff_head[3] , 
        \tx_fifo/buff_head[4] , \tx_fifo/buff_head[5] , \tx_fifo/buff_head[6] , 
        \tx_fifo/buff_head[7] , \rx_fifo/wr_index[0] , \rx_fifo/rd_index[0] , 
        \rx_fifo/length[0] , \rx_fifo/sync_wr[0] , \rx_fifo/sync_rd[0] , 
        \rx_fifo/buff_head[0] , \rx_fifo/wr_index[1] , \rx_fifo/wr_index[2] , 
        \rx_fifo/wr_index[3] , \rx_fifo/wr_index[4] , \rx_fifo/wr_index[5] , 
        \rx_fifo/wr_index[6] , \rx_fifo/wr_index[7] , \rx_fifo/rd_index[1] , 
        \rx_fifo/rd_index[2] , \rx_fifo/rd_index[3] , \rx_fifo/rd_index[4] , 
        \rx_fifo/rd_index[5] , \rx_fifo/rd_index[6] , \rx_fifo/rd_index[7] , 
        \rx_fifo/length[1] , \rx_fifo/length[2] , \rx_fifo/length[3] , 
        \rx_fifo/length[4] , \rx_fifo/length[5] , \rx_fifo/length[6] , 
        \rx_fifo/length[7] , \rx_fifo/sync_wr[1] , \rx_fifo/sync_rd[1] , 
        \i14/fifo_inst/buff[0][2] , \i14/fifo_inst/buff[0][5] , \i14/fifo_inst/buff[1][0] , 
        \i14/fifo_inst/buff[1][3] , \i14/fifo_inst/buff[1][6] , \i14/fifo_inst/buff[2][1] , 
        \i14/fifo_inst/buff[2][4] , \rx_fifo/buff_head[1] , \rx_fifo/buff_head[2] , 
        \rx_fifo/buff_head[3] , \rx_fifo/buff_head[4] , \rx_fifo/buff_head[5] , 
        \rx_fifo/buff_head[6] , \rx_fifo/buff_head[7] , \i14/fifo_inst/buff[3][3] , 
        \i14/fifo_inst/buff[3][4] , \i14/fifo_inst/buff[3][5] , \i14/fifo_inst/buff[3][6] , 
        \i14/fifo_inst/buff[3][7] , \i14/fifo_inst/buff[4][0] , \i14/fifo_inst/buff[4][1] , 
        \i14/fifo_inst/buff[4][2] , \i14/fifo_inst/buff[4][3] , \i14/fifo_inst/buff[4][4] , 
        \i14/fifo_inst/buff[4][5] , \i14/fifo_inst/buff[4][6] , \i14/fifo_inst/buff[4][7] , 
        \i14/fifo_inst/buff[5][0] , \i14/fifo_inst/buff[5][1] , \i14/fifo_inst/buff[5][2] , 
        \i14/fifo_inst/buff[5][3] , \i14/fifo_inst/buff[5][4] , \i14/fifo_inst/buff[5][5] , 
        \i14/fifo_inst/buff[5][6] , \i14/fifo_inst/buff[5][7] , \i14/fifo_inst/buff[6][0] , 
        \i14/fifo_inst/buff[6][1] , \i14/fifo_inst/buff[6][2] , \i14/fifo_inst/buff[6][3] , 
        \i14/fifo_inst/buff[6][4] , \i14/fifo_inst/buff[6][5] , \i14/fifo_inst/buff[6][6] , 
        \i14/fifo_inst/buff[6][7] , \i14/fifo_inst/buff[7][0] , \i14/fifo_inst/buff[7][1] , 
        \i14/fifo_inst/buff[7][2] , \i14/fifo_inst/buff[7][3] , \i14/fifo_inst/buff[7][4] , 
        \i14/fifo_inst/buff[7][5] , \i14/fifo_inst/buff[7][6] , \i14/fifo_inst/buff[7][7] , 
        \i14/fifo_inst/buff[8][0] , \i14/fifo_inst/buff[8][1] , \i14/fifo_inst/buff[8][2] , 
        \i14/fifo_inst/buff[8][3] , \i14/fifo_inst/buff[8][4] , \i14/fifo_inst/buff[8][5] , 
        \i14/fifo_inst/buff[8][6] , \i14/fifo_inst/buff[8][7] , \i14/fifo_inst/buff[9][0] , 
        \i14/fifo_inst/buff[9][1] , \i14/fifo_inst/buff[9][2] , \i14/fifo_inst/buff[9][3] , 
        \i14/fifo_inst/buff[9][4] , \i14/fifo_inst/buff[9][5] , \i14/fifo_inst/buff[9][6] , 
        \i14/fifo_inst/buff[9][7] , \i14/fifo_inst/buff[10][0] , \i14/fifo_inst/buff[10][1] , 
        \i14/fifo_inst/buff[10][2] , \i14/fifo_inst/buff[10][3] , \i14/fifo_inst/buff[10][4] , 
        \i14/fifo_inst/buff[10][5] , \i14/fifo_inst/buff[10][6] , \i14/fifo_inst/buff[10][7] , 
        \i14/fifo_inst/buff[11][0] , \i14/fifo_inst/buff[11][1] , \i14/fifo_inst/buff[11][2] , 
        \i14/fifo_inst/buff[11][3] , \i14/fifo_inst/buff[11][4] , \i14/fifo_inst/buff[11][5] , 
        \i14/fifo_inst/buff[11][6] , \i14/fifo_inst/buff[11][7] , \i14/fifo_inst/buff[12][0] , 
        \i14/fifo_inst/buff[12][1] , \i14/fifo_inst/buff[12][2] , \i14/fifo_inst/buff[12][3] , 
        \i14/fifo_inst/buff[12][4] , \i14/fifo_inst/buff[12][5] , \i14/fifo_inst/buff[12][6] , 
        \i14/fifo_inst/buff[12][7] , \i14/fifo_inst/buff[13][0] , \i14/fifo_inst/buff[13][1] , 
        \i14/fifo_inst/buff[13][2] , \i14/fifo_inst/buff[13][3] , \i14/fifo_inst/buff[13][4] , 
        \i14/fifo_inst/buff[13][5] , \i14/fifo_inst/buff[13][6] , \i14/fifo_inst/buff[13][7] , 
        \i14/fifo_inst/buff[14][0] , \i14/fifo_inst/buff[14][1] , \i14/fifo_inst/buff[14][2] , 
        \i14/fifo_inst/buff[14][3] , \i14/fifo_inst/buff[14][4] , \i14/fifo_inst/buff[14][5] , 
        \i14/fifo_inst/buff[14][6] , \i14/fifo_inst/buff[14][7] , \i14/fifo_inst/buff[15][0] , 
        \i14/fifo_inst/buff[15][1] , \i14/fifo_inst/buff[15][2] , \i14/fifo_inst/buff[15][3] , 
        \i14/fifo_inst/buff[15][4] , \i14/fifo_inst/buff[15][5] , \i14/fifo_inst/buff[15][6] , 
        \i14/fifo_inst/buff[15][7] , \i14/fifo_inst/buff[16][0] , \i14/fifo_inst/buff[16][1] , 
        \i14/fifo_inst/buff[16][2] , \i14/fifo_inst/buff[16][3] , \i14/fifo_inst/buff[16][4] , 
        \i14/fifo_inst/buff[16][5] , \i14/fifo_inst/buff[16][6] , \i14/fifo_inst/buff[16][7] , 
        \i14/fifo_inst/buff[17][0] , \i14/fifo_inst/buff[17][1] , \i14/fifo_inst/buff[17][2] , 
        \i14/fifo_inst/buff[17][3] , \i14/fifo_inst/buff[17][4] , \i14/fifo_inst/buff[17][5] , 
        \i14/fifo_inst/buff[17][6] , \i14/fifo_inst/buff[17][7] , \i14/fifo_inst/buff[18][0] , 
        \i14/fifo_inst/buff[18][1] , \i14/fifo_inst/buff[18][2] , \i14/fifo_inst/buff[18][3] , 
        \i14/fifo_inst/buff[18][4] , \i14/fifo_inst/buff[18][5] , \i14/fifo_inst/buff[18][6] , 
        \i14/fifo_inst/buff[18][7] , \i14/fifo_inst/buff[19][0] , \i14/fifo_inst/buff[19][1] , 
        \i14/fifo_inst/buff[19][2] , \i14/fifo_inst/buff[19][3] , \i14/fifo_inst/buff[19][4] , 
        \i14/fifo_inst/buff[19][5] , \i14/fifo_inst/buff[19][6] , \i14/fifo_inst/buff[19][7] , 
        \i14/fifo_inst/buff[20][0] , \i14/fifo_inst/buff[20][1] , \i14/fifo_inst/buff[20][2] , 
        \i14/fifo_inst/buff[20][3] , \i14/fifo_inst/buff[20][4] , \i14/fifo_inst/buff[20][5] , 
        \i14/fifo_inst/buff[20][6] , \i14/fifo_inst/buff[20][7] , \i14/fifo_inst/buff[21][0] , 
        \i14/fifo_inst/buff[21][1] , \i14/fifo_inst/buff[21][2] , \i14/fifo_inst/buff[21][3] , 
        \i14/fifo_inst/buff[21][4] , \i14/fifo_inst/buff[21][5] , \i14/fifo_inst/buff[21][6] , 
        \i14/fifo_inst/buff[21][7] , \i14/fifo_inst/buff[22][0] , \i14/fifo_inst/buff[22][1] , 
        \i14/fifo_inst/buff[22][2] , \i14/fifo_inst/buff[22][3] , \i14/fifo_inst/buff[22][4] , 
        \i14/fifo_inst/buff[22][5] , \i14/fifo_inst/buff[22][6] , \i14/fifo_inst/buff[22][7] , 
        \i14/fifo_inst/buff[23][0] , \i14/fifo_inst/buff[23][1] , \i14/fifo_inst/buff[23][2] , 
        \i14/fifo_inst/buff[23][3] , \i14/fifo_inst/buff[23][4] , \i14/fifo_inst/buff[23][5] , 
        \i14/fifo_inst/buff[23][6] , \i14/fifo_inst/buff[23][7] , \i14/fifo_inst/buff[24][0] , 
        \i14/fifo_inst/buff[24][1] , \i14/fifo_inst/buff[24][2] , \i14/fifo_inst/buff[24][3] , 
        \i14/fifo_inst/buff[24][4] , \i14/fifo_inst/buff[24][5] , \i14/fifo_inst/buff[24][6] , 
        \i14/fifo_inst/buff[24][7] , \i14/fifo_inst/buff[25][0] , \i14/fifo_inst/buff[25][1] , 
        \i14/fifo_inst/buff[25][2] , \i14/fifo_inst/buff[25][3] , \i14/fifo_inst/buff[25][4] , 
        \i14/fifo_inst/buff[25][5] , \i14/fifo_inst/buff[25][6] , \i14/fifo_inst/buff[25][7] , 
        \i14/fifo_inst/buff[26][0] , \i14/fifo_inst/buff[26][1] , \i14/fifo_inst/buff[26][2] , 
        \i14/fifo_inst/buff[26][3] , \i14/fifo_inst/buff[26][4] , \i14/fifo_inst/buff[26][5] , 
        \i14/fifo_inst/buff[26][6] , \i14/fifo_inst/buff[26][7] , \i14/fifo_inst/buff[27][0] , 
        \i14/fifo_inst/buff[27][1] , \i14/fifo_inst/buff[27][2] , \i14/fifo_inst/buff[27][3] , 
        \i14/fifo_inst/buff[27][4] , \i14/fifo_inst/buff[27][5] , \i14/fifo_inst/buff[27][6] , 
        \i14/fifo_inst/buff[27][7] , \i14/fifo_inst/buff[28][0] , \i14/fifo_inst/buff[28][1] , 
        \i14/fifo_inst/buff[28][2] , \i14/fifo_inst/buff[28][3] , \i14/fifo_inst/buff[28][4] , 
        \i14/fifo_inst/buff[28][5] , \i14/fifo_inst/buff[28][6] , \i14/fifo_inst/buff[28][7] , 
        \i14/fifo_inst/buff[29][0] , \i14/fifo_inst/buff[29][1] , \i14/fifo_inst/buff[29][2] , 
        \i14/fifo_inst/buff[29][3] , \i14/fifo_inst/buff[29][4] , \i14/fifo_inst/buff[29][5] , 
        \i14/fifo_inst/buff[29][6] , \i14/fifo_inst/buff[29][7] , \i14/fifo_inst/buff[30][0] , 
        \i14/fifo_inst/buff[30][1] , \i14/fifo_inst/buff[30][2] , \i14/fifo_inst/buff[30][3] , 
        \i14/fifo_inst/buff[30][4] , \i14/fifo_inst/buff[30][5] , \i14/fifo_inst/buff[30][6] , 
        \i14/fifo_inst/buff[30][7] , \i14/fifo_inst/buff[31][0] , \i14/fifo_inst/buff[31][1] , 
        \i14/fifo_inst/buff[31][2] , \i14/fifo_inst/buff[31][3] , \i14/fifo_inst/buff[31][4] , 
        \i14/fifo_inst/buff[31][5] , \i14/fifo_inst/buff[31][6] , \i14/fifo_inst/buff[31][7] , 
        \i14/fifo_inst/buff[32][0] , \i14/fifo_inst/buff[32][1] , \i14/fifo_inst/buff[32][2] , 
        \i14/fifo_inst/buff[32][3] , \i14/fifo_inst/buff[32][4] , \i14/fifo_inst/buff[32][5] , 
        \i14/fifo_inst/buff[32][6] , \i14/fifo_inst/buff[32][7] , \i14/fifo_inst/buff[33][0] , 
        \i14/fifo_inst/buff[33][1] , \i14/fifo_inst/buff[33][2] , \i14/fifo_inst/buff[33][3] , 
        \i14/fifo_inst/buff[33][4] , \i14/fifo_inst/buff[33][5] , \i14/fifo_inst/buff[33][6] , 
        \i14/fifo_inst/buff[33][7] , \i14/fifo_inst/buff[34][0] , \i14/fifo_inst/buff[34][1] , 
        \i14/fifo_inst/buff[34][2] , \i14/fifo_inst/buff[34][3] , \i14/fifo_inst/buff[34][4] , 
        \i14/fifo_inst/buff[34][5] , \i14/fifo_inst/buff[34][6] , \i14/fifo_inst/buff[34][7] , 
        \i14/fifo_inst/buff[35][0] , \i14/fifo_inst/buff[35][1] , \i14/fifo_inst/buff[35][2] , 
        \i14/fifo_inst/buff[35][3] , \i14/fifo_inst/buff[35][4] , \i14/fifo_inst/buff[35][5] , 
        \i14/fifo_inst/buff[35][6] , \i14/fifo_inst/buff[35][7] , \i14/fifo_inst/buff[36][0] , 
        \i14/fifo_inst/buff[36][1] , \i14/fifo_inst/buff[36][2] , \i14/fifo_inst/buff[36][3] , 
        \i14/fifo_inst/buff[36][4] , \i14/fifo_inst/buff[36][5] , \i14/fifo_inst/buff[36][6] , 
        \i14/fifo_inst/buff[36][7] , \i14/fifo_inst/buff[37][0] , \i14/fifo_inst/buff[37][1] , 
        \i14/fifo_inst/buff[37][2] , \i14/fifo_inst/buff[37][3] , \i14/fifo_inst/buff[37][4] , 
        \i14/fifo_inst/buff[37][5] , \i14/fifo_inst/buff[37][6] , \i14/fifo_inst/buff[37][7] , 
        \i14/fifo_inst/buff[38][0] , \i14/fifo_inst/buff[38][1] , \i14/fifo_inst/buff[38][2] , 
        \i14/fifo_inst/buff[38][3] , \i14/fifo_inst/buff[38][4] , \i14/fifo_inst/buff[38][5] , 
        \i14/fifo_inst/buff[38][6] , \i14/fifo_inst/buff[38][7] , \i14/fifo_inst/buff[39][0] , 
        \i14/fifo_inst/buff[39][1] , \i14/fifo_inst/buff[39][2] , \i14/fifo_inst/buff[39][3] , 
        \i14/fifo_inst/buff[39][4] , \i14/fifo_inst/buff[39][5] , \i14/fifo_inst/buff[39][6] , 
        \i14/fifo_inst/buff[39][7] , \i14/fifo_inst/buff[40][0] , \i14/fifo_inst/buff[40][1] , 
        \i14/fifo_inst/buff[40][2] , \i14/fifo_inst/buff[40][3] , \i14/fifo_inst/buff[40][4] , 
        \i14/fifo_inst/buff[40][5] , \i14/fifo_inst/buff[40][6] , \i14/fifo_inst/buff[40][7] , 
        \i14/fifo_inst/buff[41][0] , \i14/fifo_inst/buff[41][1] , \i14/fifo_inst/buff[41][2] , 
        \i14/fifo_inst/buff[41][3] , \i14/fifo_inst/buff[41][4] , \i14/fifo_inst/buff[41][5] , 
        \i14/fifo_inst/buff[41][6] , \i14/fifo_inst/buff[41][7] , \i14/fifo_inst/buff[42][0] , 
        \i14/fifo_inst/buff[42][1] , \i14/fifo_inst/buff[42][2] , \i14/fifo_inst/buff[42][3] , 
        \i14/fifo_inst/buff[42][4] , \i14/fifo_inst/buff[42][5] , \i14/fifo_inst/buff[42][6] , 
        \i14/fifo_inst/buff[42][7] , \i14/fifo_inst/buff[43][0] , \i14/fifo_inst/buff[43][1] , 
        \i14/fifo_inst/buff[43][2] , \i14/fifo_inst/buff[43][3] , \i14/fifo_inst/buff[43][4] , 
        \i14/fifo_inst/buff[43][5] , \i14/fifo_inst/buff[43][6] , \i14/fifo_inst/buff[43][7] , 
        \i14/fifo_inst/buff[44][0] , \i14/fifo_inst/buff[44][1] , \i14/fifo_inst/buff[44][2] , 
        \i14/fifo_inst/buff[44][3] , \i14/fifo_inst/buff[44][4] , \i14/fifo_inst/buff[44][5] , 
        \i14/fifo_inst/buff[44][6] , \i14/fifo_inst/buff[44][7] , \i14/fifo_inst/buff[45][0] , 
        \i14/fifo_inst/buff[45][1] , \i14/fifo_inst/buff[45][2] , \i14/fifo_inst/buff[45][3] , 
        \i14/fifo_inst/buff[45][4] , \i14/fifo_inst/buff[45][5] , \i14/fifo_inst/buff[45][6] , 
        \i14/fifo_inst/buff[45][7] , \i14/fifo_inst/buff[46][0] , \i14/fifo_inst/buff[46][1] , 
        \i14/fifo_inst/buff[46][2] , \i14/fifo_inst/buff[46][3] , \i14/fifo_inst/buff[46][4] , 
        \i14/fifo_inst/buff[46][5] , \i14/fifo_inst/buff[46][6] , \i14/fifo_inst/buff[46][7] , 
        \i14/fifo_inst/buff[47][0] , \i14/fifo_inst/buff[47][1] , \i14/fifo_inst/buff[47][2] , 
        \i14/fifo_inst/buff[47][3] , \i14/fifo_inst/buff[47][4] , \i14/fifo_inst/buff[47][5] , 
        \i14/fifo_inst/buff[47][6] , \i14/fifo_inst/buff[47][7] , \i14/fifo_inst/buff[48][0] , 
        \i14/fifo_inst/buff[48][1] , \i14/fifo_inst/buff[48][2] , \i14/fifo_inst/buff[48][3] , 
        \i14/fifo_inst/buff[48][4] , \i14/fifo_inst/buff[48][5] , \i14/fifo_inst/buff[48][6] , 
        \i14/fifo_inst/buff[48][7] , \i14/fifo_inst/buff[49][0] , \i14/fifo_inst/buff[49][1] , 
        \i14/fifo_inst/buff[49][2] , \i14/fifo_inst/buff[49][3] , \i14/fifo_inst/buff[49][4] , 
        \i14/fifo_inst/buff[49][5] , \i14/fifo_inst/buff[49][6] , \i14/fifo_inst/buff[49][7] , 
        \i14/fifo_inst/buff[50][0] , \i14/fifo_inst/buff[50][1] , \i14/fifo_inst/buff[50][2] , 
        \i14/fifo_inst/buff[50][3] , \i14/fifo_inst/buff[50][4] , \i14/fifo_inst/buff[50][5] , 
        \i14/fifo_inst/buff[50][6] , \i14/fifo_inst/buff[50][7] , \i14/fifo_inst/buff[51][0] , 
        \i14/fifo_inst/buff[51][1] , \i14/fifo_inst/buff[51][2] , \i14/fifo_inst/buff[51][3] , 
        \i14/fifo_inst/buff[51][4] , \i14/fifo_inst/buff[51][5] , \i14/fifo_inst/buff[51][6] , 
        \i14/fifo_inst/buff[51][7] , \i14/fifo_inst/buff[52][0] , \i14/fifo_inst/buff[52][1] , 
        \i14/fifo_inst/buff[52][2] , \i14/fifo_inst/buff[52][3] , \i14/fifo_inst/buff[52][4] , 
        \i14/fifo_inst/buff[52][5] , \i14/fifo_inst/buff[52][6] , \i14/fifo_inst/buff[52][7] , 
        \i14/fifo_inst/buff[53][0] , \i14/fifo_inst/buff[53][1] , \i14/fifo_inst/buff[53][2] , 
        \i14/fifo_inst/buff[53][3] , \i14/fifo_inst/buff[53][4] , \i14/fifo_inst/buff[53][5] , 
        \i14/fifo_inst/buff[53][6] , \i14/fifo_inst/buff[53][7] , \i14/fifo_inst/buff[54][0] , 
        \i14/fifo_inst/buff[54][1] , \i14/fifo_inst/buff[54][2] , \i14/fifo_inst/buff[54][3] , 
        \i14/fifo_inst/buff[54][4] , \i14/fifo_inst/buff[54][5] , \i14/fifo_inst/buff[54][6] , 
        \i14/fifo_inst/buff[54][7] , \i14/fifo_inst/buff[55][0] , \i14/fifo_inst/buff[55][1] , 
        \i14/fifo_inst/buff[55][2] , \i14/fifo_inst/buff[55][3] , \i14/fifo_inst/buff[55][4] , 
        \i14/fifo_inst/buff[55][5] , \i14/fifo_inst/buff[55][6] , \i14/fifo_inst/buff[55][7] , 
        \i14/fifo_inst/buff[56][0] , \i14/fifo_inst/buff[56][1] , \i14/fifo_inst/buff[56][2] , 
        \i14/fifo_inst/buff[56][3] , \i14/fifo_inst/buff[56][4] , \i14/fifo_inst/buff[56][5] , 
        \i14/fifo_inst/buff[56][6] , \i14/fifo_inst/buff[56][7] , \i14/fifo_inst/buff[57][0] , 
        \i14/fifo_inst/buff[57][1] , \i14/fifo_inst/buff[57][2] , \i14/fifo_inst/buff[57][3] , 
        \i14/fifo_inst/buff[57][4] , \i14/fifo_inst/buff[57][5] , \i14/fifo_inst/buff[57][6] , 
        \i14/fifo_inst/buff[57][7] , \i14/fifo_inst/buff[58][0] , \i14/fifo_inst/buff[58][1] , 
        \i14/fifo_inst/buff[58][2] , \i14/fifo_inst/buff[58][3] , \i14/fifo_inst/buff[58][4] , 
        \i14/fifo_inst/buff[58][5] , \i14/fifo_inst/buff[58][6] , \i14/fifo_inst/buff[58][7] , 
        \i14/fifo_inst/buff[59][0] , \i14/fifo_inst/buff[59][1] , \i14/fifo_inst/buff[59][2] , 
        \i14/fifo_inst/buff[59][3] , \i14/fifo_inst/buff[59][4] , \i14/fifo_inst/buff[59][5] , 
        \i14/fifo_inst/buff[59][6] , \i14/fifo_inst/buff[59][7] , \i14/fifo_inst/buff[60][0] , 
        \i14/fifo_inst/buff[60][1] , \i14/fifo_inst/buff[60][2] , \i14/fifo_inst/buff[60][3] , 
        \i14/fifo_inst/buff[60][4] , \i14/fifo_inst/buff[60][5] , \i14/fifo_inst/buff[60][6] , 
        \i14/fifo_inst/buff[60][7] , \i14/fifo_inst/buff[61][0] , \i14/fifo_inst/buff[61][1] , 
        \i14/fifo_inst/buff[61][2] , \i14/fifo_inst/buff[61][3] , \i14/fifo_inst/buff[61][4] , 
        \i14/fifo_inst/buff[61][5] , \i14/fifo_inst/buff[61][6] , \i14/fifo_inst/buff[61][7] , 
        \i14/fifo_inst/buff[62][0] , \i14/fifo_inst/buff[62][1] , \i14/fifo_inst/buff[62][2] , 
        \i14/fifo_inst/buff[62][3] , \i14/fifo_inst/buff[62][4] , \i14/fifo_inst/buff[62][5] , 
        \i14/fifo_inst/buff[62][6] , \i14/fifo_inst/buff[62][7] , \i14/fifo_inst/buff[63][0] , 
        \i14/fifo_inst/buff[63][1] , \i14/fifo_inst/buff[63][2] , \i14/fifo_inst/buff[63][3] , 
        \i14/fifo_inst/buff[63][4] , \i14/fifo_inst/buff[63][5] , \i14/fifo_inst/buff[63][6] , 
        \i14/fifo_inst/buff[63][7] , \i14/fifo_inst/buff[64][0] , \i14/fifo_inst/buff[64][1] , 
        \i14/fifo_inst/buff[64][2] , \i14/fifo_inst/buff[64][3] , \i14/fifo_inst/buff[64][4] , 
        \i14/fifo_inst/buff[64][5] , \i14/fifo_inst/buff[64][6] , \i14/fifo_inst/buff[64][7] , 
        \i14/fifo_inst/buff[65][0] , \i14/fifo_inst/buff[65][1] , \i14/fifo_inst/buff[65][2] , 
        \i14/fifo_inst/buff[65][3] , \i14/fifo_inst/buff[65][4] , \i14/fifo_inst/buff[65][5] , 
        \i14/fifo_inst/buff[65][6] , \i14/fifo_inst/buff[65][7] , \i14/fifo_inst/buff[66][0] , 
        \i14/fifo_inst/buff[66][1] , \i14/fifo_inst/buff[66][2] , \i14/fifo_inst/buff[66][3] , 
        \i14/fifo_inst/buff[66][4] , \i14/fifo_inst/buff[66][5] , \i14/fifo_inst/buff[66][6] , 
        \i14/fifo_inst/buff[66][7] , \i14/fifo_inst/buff[67][0] , \i14/fifo_inst/buff[67][1] , 
        \i14/fifo_inst/buff[67][2] , \i14/fifo_inst/buff[67][3] , \i14/fifo_inst/buff[67][4] , 
        \i14/fifo_inst/buff[67][5] , \i14/fifo_inst/buff[67][6] , \i14/fifo_inst/buff[67][7] , 
        \i14/fifo_inst/buff[68][0] , \i14/fifo_inst/buff[68][1] , \i14/fifo_inst/buff[68][2] , 
        \i14/fifo_inst/buff[68][3] , \i14/fifo_inst/buff[68][4] , \i14/fifo_inst/buff[68][5] , 
        \i14/fifo_inst/buff[68][6] , \i14/fifo_inst/buff[68][7] , \i14/fifo_inst/buff[69][0] , 
        \i14/fifo_inst/buff[69][1] , \i14/fifo_inst/buff[69][2] , \i14/fifo_inst/buff[69][3] , 
        \i14/fifo_inst/buff[69][4] , \i14/fifo_inst/buff[69][5] , \i14/fifo_inst/buff[69][6] , 
        \i14/fifo_inst/buff[69][7] , \i14/fifo_inst/buff[70][0] , \i14/fifo_inst/buff[70][1] , 
        \i14/fifo_inst/buff[70][2] , \i14/fifo_inst/buff[70][3] , \i14/fifo_inst/buff[70][4] , 
        \i14/fifo_inst/buff[70][5] , \i14/fifo_inst/buff[70][6] , \i14/fifo_inst/buff[70][7] , 
        \i14/fifo_inst/buff[71][0] , \i14/fifo_inst/buff[71][1] , \i14/fifo_inst/buff[71][2] , 
        \i14/fifo_inst/buff[71][3] , \i14/fifo_inst/buff[71][4] , \i14/fifo_inst/buff[71][5] , 
        \i14/fifo_inst/buff[71][6] , \i14/fifo_inst/buff[71][7] , \i14/fifo_inst/buff[72][0] , 
        \i14/fifo_inst/buff[72][1] , \i14/fifo_inst/buff[72][2] , \i14/fifo_inst/buff[72][3] , 
        \i14/fifo_inst/buff[72][4] , \i14/fifo_inst/buff[72][5] , \i14/fifo_inst/buff[72][6] , 
        \i14/fifo_inst/buff[72][7] , \i14/fifo_inst/buff[73][0] , \i14/fifo_inst/buff[73][1] , 
        \i14/fifo_inst/buff[73][2] , \i14/fifo_inst/buff[73][3] , \i14/fifo_inst/buff[73][4] , 
        \i14/fifo_inst/buff[73][5] , \i14/fifo_inst/buff[73][6] , \i14/fifo_inst/buff[73][7] , 
        \i14/fifo_inst/buff[74][0] , \i14/fifo_inst/buff[74][1] , \i14/fifo_inst/buff[74][2] , 
        \i14/fifo_inst/buff[74][3] , \i14/fifo_inst/buff[74][4] , \i14/fifo_inst/buff[74][5] , 
        \i14/fifo_inst/buff[74][6] , \i14/fifo_inst/buff[74][7] , \i14/fifo_inst/buff[75][0] , 
        \i14/fifo_inst/buff[75][1] , \i14/fifo_inst/buff[75][2] , \i14/fifo_inst/buff[75][3] , 
        \i14/fifo_inst/buff[75][4] , \i14/fifo_inst/buff[75][5] , \i14/fifo_inst/buff[75][6] , 
        \i14/fifo_inst/buff[75][7] , \i14/fifo_inst/buff[76][0] , \i14/fifo_inst/buff[76][1] , 
        \i14/fifo_inst/buff[76][2] , \i14/fifo_inst/buff[76][3] , \i14/fifo_inst/buff[76][4] , 
        \i14/fifo_inst/buff[76][5] , \i14/fifo_inst/buff[76][6] , \i14/fifo_inst/buff[76][7] , 
        \i14/fifo_inst/buff[77][0] , \i14/fifo_inst/buff[77][1] , \i14/fifo_inst/buff[77][2] , 
        \i14/fifo_inst/buff[77][3] , \i14/fifo_inst/buff[77][4] , \i14/fifo_inst/buff[77][5] , 
        \i14/fifo_inst/buff[77][6] , \i14/fifo_inst/buff[77][7] , \i14/fifo_inst/buff[78][0] , 
        \i14/fifo_inst/buff[78][1] , \i14/fifo_inst/buff[78][2] , \i14/fifo_inst/buff[78][3] , 
        \i14/fifo_inst/buff[78][4] , \i14/fifo_inst/buff[78][5] , \i14/fifo_inst/buff[78][6] , 
        \i14/fifo_inst/buff[78][7] , \i14/fifo_inst/buff[79][0] , \i14/fifo_inst/buff[79][1] , 
        \i14/fifo_inst/buff[79][2] , \i14/fifo_inst/buff[79][3] , \i14/fifo_inst/buff[79][4] , 
        \i14/fifo_inst/buff[79][5] , \i14/fifo_inst/buff[79][6] , \i14/fifo_inst/buff[79][7] , 
        \i14/fifo_inst/buff[80][0] , \i14/fifo_inst/buff[80][1] , \i14/fifo_inst/buff[80][2] , 
        \i14/fifo_inst/buff[80][3] , \i14/fifo_inst/buff[80][4] , \i14/fifo_inst/buff[80][5] , 
        \i14/fifo_inst/buff[80][6] , \i14/fifo_inst/buff[80][7] , \i14/fifo_inst/buff[81][0] , 
        \i14/fifo_inst/buff[81][1] , \i14/fifo_inst/buff[81][2] , \i14/fifo_inst/buff[81][3] , 
        \i14/fifo_inst/buff[81][4] , \i14/fifo_inst/buff[81][5] , \i14/fifo_inst/buff[81][6] , 
        \i14/fifo_inst/buff[81][7] , \i14/fifo_inst/buff[82][0] , \i14/fifo_inst/buff[82][1] , 
        \i14/fifo_inst/buff[82][2] , \i14/fifo_inst/buff[82][3] , \i14/fifo_inst/buff[82][4] , 
        \i14/fifo_inst/buff[82][5] , \i14/fifo_inst/buff[82][6] , \i14/fifo_inst/buff[82][7] , 
        \i14/fifo_inst/buff[83][0] , \i14/fifo_inst/buff[83][1] , \i14/fifo_inst/buff[83][2] , 
        \i14/fifo_inst/buff[83][3] , \i14/fifo_inst/buff[83][4] , \i14/fifo_inst/buff[83][5] , 
        \i14/fifo_inst/buff[83][6] , \i14/fifo_inst/buff[83][7] , \i14/fifo_inst/buff[84][0] , 
        \i14/fifo_inst/buff[84][1] , \i14/fifo_inst/buff[84][2] , \i14/fifo_inst/buff[84][3] , 
        \i14/fifo_inst/buff[84][4] , \i14/fifo_inst/buff[84][5] , \i14/fifo_inst/buff[84][6] , 
        \i14/fifo_inst/buff[84][7] , \i14/fifo_inst/buff[85][0] , \i14/fifo_inst/buff[85][1] , 
        \i14/fifo_inst/buff[85][2] , \i14/fifo_inst/buff[85][3] , \i14/fifo_inst/buff[85][4] , 
        \i14/fifo_inst/buff[85][5] , \i14/fifo_inst/buff[85][6] , \i14/fifo_inst/buff[85][7] , 
        \i14/fifo_inst/buff[86][0] , \i14/fifo_inst/buff[86][1] , \i14/fifo_inst/buff[86][2] , 
        \i14/fifo_inst/buff[86][3] , \i14/fifo_inst/buff[86][4] , \i14/fifo_inst/buff[86][5] , 
        \i14/fifo_inst/buff[86][6] , \i14/fifo_inst/buff[86][7] , \i14/fifo_inst/buff[87][0] , 
        \i14/fifo_inst/buff[87][1] , \i14/fifo_inst/buff[87][2] , \i14/fifo_inst/buff[87][3] , 
        \i14/fifo_inst/buff[87][4] , \i14/fifo_inst/buff[87][5] , \i14/fifo_inst/buff[87][6] , 
        \i14/fifo_inst/buff[87][7] , \i14/fifo_inst/buff[88][0] , \i14/fifo_inst/buff[88][1] , 
        \i14/fifo_inst/buff[88][2] , \i14/fifo_inst/buff[88][3] , \i14/fifo_inst/buff[88][4] , 
        \i14/fifo_inst/buff[88][5] , \i14/fifo_inst/buff[88][6] , \i14/fifo_inst/buff[88][7] , 
        \i14/fifo_inst/buff[89][0] , \i14/fifo_inst/buff[89][1] , \i14/fifo_inst/buff[89][2] , 
        \i14/fifo_inst/buff[89][3] , \i14/fifo_inst/buff[89][4] , \i14/fifo_inst/buff[89][5] , 
        \i14/fifo_inst/buff[89][6] , \i14/fifo_inst/buff[89][7] , \i14/fifo_inst/buff[90][0] , 
        \i14/fifo_inst/buff[90][1] , \i14/fifo_inst/buff[90][2] , \i14/fifo_inst/buff[90][3] , 
        \i14/fifo_inst/buff[90][4] , \i14/fifo_inst/buff[90][5] , \i14/fifo_inst/buff[90][6] , 
        \i14/fifo_inst/buff[90][7] , \i14/fifo_inst/buff[91][0] , \i14/fifo_inst/buff[91][1] , 
        \i14/fifo_inst/buff[91][2] , \i14/fifo_inst/buff[91][3] , \i14/fifo_inst/buff[91][4] , 
        \i14/fifo_inst/buff[91][5] , \i14/fifo_inst/buff[91][6] , \i14/fifo_inst/buff[91][7] , 
        \i14/fifo_inst/buff[92][0] , \i14/fifo_inst/buff[92][1] , \i14/fifo_inst/buff[92][2] , 
        \i14/fifo_inst/buff[92][3] , \i14/fifo_inst/buff[92][4] , \i14/fifo_inst/buff[92][5] , 
        \i14/fifo_inst/buff[92][6] , \i14/fifo_inst/buff[92][7] , \i14/fifo_inst/buff[93][0] , 
        \i14/fifo_inst/buff[93][1] , \i14/fifo_inst/buff[93][2] , \i14/fifo_inst/buff[93][3] , 
        \i14/fifo_inst/buff[93][4] , \i14/fifo_inst/buff[93][5] , \i14/fifo_inst/buff[93][6] , 
        \i14/fifo_inst/buff[93][7] , \i14/fifo_inst/buff[94][0] , \i14/fifo_inst/buff[94][1] , 
        \i14/fifo_inst/buff[94][2] , \i14/fifo_inst/buff[94][3] , \i14/fifo_inst/buff[94][4] , 
        \i14/fifo_inst/buff[94][5] , \i14/fifo_inst/buff[94][6] , \i14/fifo_inst/buff[94][7] , 
        \i14/fifo_inst/buff[95][0] , \i14/fifo_inst/buff[95][1] , \i14/fifo_inst/buff[95][2] , 
        \i14/fifo_inst/buff[95][3] , \i14/fifo_inst/buff[95][4] , \i14/fifo_inst/buff[95][5] , 
        \i14/fifo_inst/buff[95][6] , \i14/fifo_inst/buff[95][7] , \i14/fifo_inst/buff[96][0] , 
        \i14/fifo_inst/buff[96][1] , \i14/fifo_inst/buff[96][2] , \i14/fifo_inst/buff[96][3] , 
        \i14/fifo_inst/buff[96][4] , \i14/fifo_inst/buff[96][5] , \i14/fifo_inst/buff[96][6] , 
        \i14/fifo_inst/buff[96][7] , \i14/fifo_inst/buff[97][0] , \i14/fifo_inst/buff[97][1] , 
        \i14/fifo_inst/buff[97][2] , \i14/fifo_inst/buff[97][3] , \i14/fifo_inst/buff[97][4] , 
        \i14/fifo_inst/buff[97][5] , \i14/fifo_inst/buff[97][6] , \i14/fifo_inst/buff[97][7] , 
        \i14/fifo_inst/buff[98][0] , \i14/fifo_inst/buff[98][1] , \i14/fifo_inst/buff[98][2] , 
        \i14/fifo_inst/buff[98][3] , \i14/fifo_inst/buff[98][4] , \i14/fifo_inst/buff[98][5] , 
        \i14/fifo_inst/buff[98][6] , \i14/fifo_inst/buff[98][7] , \i14/fifo_inst/buff[99][0] , 
        \i14/fifo_inst/buff[99][1] , \i14/fifo_inst/buff[99][2] , \i14/fifo_inst/buff[99][3] , 
        \i14/fifo_inst/buff[99][4] , \i14/fifo_inst/buff[99][5] , \i14/fifo_inst/buff[99][6] , 
        \i14/fifo_inst/buff[99][7] , \i14/fifo_inst/buff[100][0] , \i14/fifo_inst/buff[100][1] , 
        \i14/fifo_inst/buff[100][2] , \i14/fifo_inst/buff[100][3] , \i14/fifo_inst/buff[100][4] , 
        \i14/fifo_inst/buff[100][5] , \i14/fifo_inst/buff[100][6] , \i14/fifo_inst/buff[100][7] , 
        \i14/fifo_inst/buff[101][0] , \i14/fifo_inst/buff[101][1] , \i14/fifo_inst/buff[101][2] , 
        \i14/fifo_inst/buff[101][3] , \i14/fifo_inst/buff[101][4] , \i14/fifo_inst/buff[101][5] , 
        \i14/fifo_inst/buff[101][6] , \i14/fifo_inst/buff[101][7] , \i14/fifo_inst/buff[102][0] , 
        \i14/fifo_inst/buff[102][1] , \i14/fifo_inst/buff[102][2] , \i14/fifo_inst/buff[102][3] , 
        \i14/fifo_inst/buff[102][4] , \i14/fifo_inst/buff[102][5] , \i14/fifo_inst/buff[102][6] , 
        \i14/fifo_inst/buff[102][7] , \i14/fifo_inst/buff[103][0] , \i14/fifo_inst/buff[103][1] , 
        \i14/fifo_inst/buff[103][2] , \i14/fifo_inst/buff[103][3] , \i14/fifo_inst/buff[103][4] , 
        \i14/fifo_inst/buff[103][5] , \i14/fifo_inst/buff[103][6] , \i14/fifo_inst/buff[103][7] , 
        \i14/fifo_inst/buff[104][0] , \i14/fifo_inst/buff[104][1] , \i14/fifo_inst/buff[104][2] , 
        \i14/fifo_inst/buff[104][3] , \i14/fifo_inst/buff[104][4] , \i14/fifo_inst/buff[104][5] , 
        \i14/fifo_inst/buff[104][6] , \i14/fifo_inst/buff[104][7] , \i14/fifo_inst/buff[105][0] , 
        \i14/fifo_inst/buff[105][1] , \i14/fifo_inst/buff[105][2] , \i14/fifo_inst/buff[105][3] , 
        \i14/fifo_inst/buff[105][4] , \i14/fifo_inst/buff[105][5] , \i14/fifo_inst/buff[105][6] , 
        \i14/fifo_inst/buff[105][7] , \i14/fifo_inst/buff[106][0] , \i14/fifo_inst/buff[106][1] , 
        \i14/fifo_inst/buff[106][2] , \i14/fifo_inst/buff[106][3] , \i14/fifo_inst/buff[106][4] , 
        \i14/fifo_inst/buff[106][5] , \i14/fifo_inst/buff[106][6] , \i14/fifo_inst/buff[106][7] , 
        \i14/fifo_inst/buff[107][0] , \i14/fifo_inst/buff[107][1] , \i14/fifo_inst/buff[107][2] , 
        \i14/fifo_inst/buff[107][3] , \i14/fifo_inst/buff[107][4] , \i14/fifo_inst/buff[107][5] , 
        \i14/fifo_inst/buff[107][6] , \i14/fifo_inst/buff[107][7] , \i14/fifo_inst/buff[108][0] , 
        \i14/fifo_inst/buff[108][1] , \i14/fifo_inst/buff[108][2] , \i14/fifo_inst/buff[108][3] , 
        \i14/fifo_inst/buff[108][4] , \i14/fifo_inst/buff[108][5] , \i14/fifo_inst/buff[108][6] , 
        \i14/fifo_inst/buff[108][7] , \i14/fifo_inst/buff[109][0] , \i14/fifo_inst/buff[109][1] , 
        \i14/fifo_inst/buff[109][2] , \i14/fifo_inst/buff[109][3] , \i14/fifo_inst/buff[109][4] , 
        \i14/fifo_inst/buff[109][5] , \i14/fifo_inst/buff[109][6] , \i14/fifo_inst/buff[109][7] , 
        \i14/fifo_inst/buff[110][0] , \i14/fifo_inst/buff[110][1] , \i14/fifo_inst/buff[110][2] , 
        \i14/fifo_inst/buff[110][3] , \i14/fifo_inst/buff[110][4] , \i14/fifo_inst/buff[110][5] , 
        \i14/fifo_inst/buff[110][6] , \i14/fifo_inst/buff[110][7] , \i14/fifo_inst/buff[111][0] , 
        \i14/fifo_inst/buff[111][1] , \i14/fifo_inst/buff[111][2] , \i14/fifo_inst/buff[111][3] , 
        \i14/fifo_inst/buff[111][4] , \i14/fifo_inst/buff[111][5] , \i14/fifo_inst/buff[111][6] , 
        \i14/fifo_inst/buff[111][7] , \i14/fifo_inst/buff[112][0] , \i14/fifo_inst/buff[112][1] , 
        \i14/fifo_inst/buff[112][2] , \i14/fifo_inst/buff[112][3] , \i14/fifo_inst/buff[112][4] , 
        \i14/fifo_inst/buff[112][5] , \i14/fifo_inst/buff[112][6] , \i14/fifo_inst/buff[112][7] , 
        \i14/fifo_inst/buff[113][0] , \i14/fifo_inst/buff[113][1] , \i14/fifo_inst/buff[113][2] , 
        \i14/fifo_inst/buff[113][3] , \i14/fifo_inst/buff[113][4] , \i14/fifo_inst/buff[113][5] , 
        \i14/fifo_inst/buff[113][6] , \i14/fifo_inst/buff[113][7] , \i14/fifo_inst/buff[114][0] , 
        \i14/fifo_inst/buff[114][1] , \i14/fifo_inst/buff[114][2] , \i14/fifo_inst/buff[114][3] , 
        \i14/fifo_inst/buff[114][4] , \i14/fifo_inst/buff[114][5] , \i14/fifo_inst/buff[114][6] , 
        \i14/fifo_inst/buff[114][7] , \i14/fifo_inst/buff[115][0] , \i14/fifo_inst/buff[115][1] , 
        \i14/fifo_inst/buff[115][2] , \i14/fifo_inst/buff[115][3] , \i14/fifo_inst/buff[115][4] , 
        \i14/fifo_inst/buff[115][5] , \i14/fifo_inst/buff[115][6] , \i14/fifo_inst/buff[115][7] , 
        \i14/fifo_inst/buff[116][0] , \i14/fifo_inst/buff[116][1] , \i14/fifo_inst/buff[116][2] , 
        \i14/fifo_inst/buff[116][3] , \i14/fifo_inst/buff[116][4] , \i14/fifo_inst/buff[116][5] , 
        \i14/fifo_inst/buff[116][6] , \i14/fifo_inst/buff[116][7] , \i14/fifo_inst/buff[117][0] , 
        \i14/fifo_inst/buff[117][1] , \i14/fifo_inst/buff[117][2] , \i14/fifo_inst/buff[117][3] , 
        \i14/fifo_inst/buff[117][4] , \i14/fifo_inst/buff[117][5] , \i14/fifo_inst/buff[117][6] , 
        \i14/fifo_inst/buff[117][7] , \i14/fifo_inst/buff[118][0] , \i14/fifo_inst/buff[118][1] , 
        \i14/fifo_inst/buff[118][2] , \i14/fifo_inst/buff[118][3] , \i14/fifo_inst/buff[118][4] , 
        \i14/fifo_inst/buff[118][5] , \i14/fifo_inst/buff[118][6] , \i14/fifo_inst/buff[118][7] , 
        \i14/fifo_inst/buff[119][0] , \i14/fifo_inst/buff[119][1] , \i14/fifo_inst/buff[119][2] , 
        \i14/fifo_inst/buff[119][3] , \i14/fifo_inst/buff[119][4] , \i14/fifo_inst/buff[119][5] , 
        \i14/fifo_inst/buff[119][6] , \i14/fifo_inst/buff[119][7] , \i14/fifo_inst/buff[120][0] , 
        \i14/fifo_inst/buff[120][1] , \i14/fifo_inst/buff[120][2] , \i14/fifo_inst/buff[120][3] , 
        \i14/fifo_inst/buff[120][4] , \i14/fifo_inst/buff[120][5] , \i14/fifo_inst/buff[120][6] , 
        \i14/fifo_inst/buff[120][7] , \i14/fifo_inst/buff[121][0] , \i14/fifo_inst/buff[121][1] , 
        \i14/fifo_inst/buff[121][2] , \i14/fifo_inst/buff[121][3] , \i14/fifo_inst/buff[121][4] , 
        \i14/fifo_inst/buff[121][5] , \i14/fifo_inst/buff[121][6] , \i14/fifo_inst/buff[121][7] , 
        \i14/fifo_inst/buff[122][0] , \i14/fifo_inst/buff[122][1] , \i14/fifo_inst/buff[122][2] , 
        \i14/fifo_inst/buff[122][3] , \i14/fifo_inst/buff[122][4] , \i14/fifo_inst/buff[122][5] , 
        \i14/fifo_inst/buff[122][6] , \i14/fifo_inst/buff[122][7] , \i14/fifo_inst/buff[123][0] , 
        \i14/fifo_inst/buff[123][1] , \i14/fifo_inst/buff[123][2] , \i14/fifo_inst/buff[123][3] , 
        \i14/fifo_inst/buff[123][4] , \i14/fifo_inst/buff[123][5] , \i14/fifo_inst/buff[123][6] , 
        \i14/fifo_inst/buff[123][7] , \i14/fifo_inst/buff[124][0] , \i14/fifo_inst/buff[124][1] , 
        \i14/fifo_inst/buff[124][2] , \i14/fifo_inst/buff[124][3] , \i14/fifo_inst/buff[124][4] , 
        \i14/fifo_inst/buff[124][5] , \i14/fifo_inst/buff[124][6] , \i14/fifo_inst/buff[124][7] , 
        \i14/fifo_inst/buff[125][0] , \i14/fifo_inst/buff[125][1] , \i14/fifo_inst/buff[125][2] , 
        \i14/fifo_inst/buff[125][3] , \i14/fifo_inst/buff[125][4] , \i14/fifo_inst/buff[125][5] , 
        \i14/fifo_inst/buff[125][6] , \i14/fifo_inst/buff[125][7] , \i14/fifo_inst/buff[126][0] , 
        \i14/fifo_inst/buff[126][1] , \i14/fifo_inst/buff[126][2] , \i14/fifo_inst/buff[126][3] , 
        \i14/fifo_inst/buff[126][4] , \i14/fifo_inst/buff[126][5] , \i14/fifo_inst/buff[126][6] , 
        \i14/fifo_inst/buff[126][7] , \i14/fifo_inst/buff[127][0] , \i14/fifo_inst/buff[127][1] , 
        \i14/fifo_inst/buff[127][2] , \i14/fifo_inst/buff[127][3] , \i14/fifo_inst/buff[127][4] , 
        \i14/fifo_inst/buff[127][5] , \i14/fifo_inst/buff[127][6] , \i14/fifo_inst/buff[127][7] , 
        \i15/tx_fifo/buff[0][0] , \i15/tx_fifo/buff[0][1] , \i15/tx_fifo/buff[0][2] , 
        \i15/tx_fifo/buff[0][3] , \i15/tx_fifo/buff[0][4] , \i15/tx_fifo/buff[0][5] , 
        \i15/tx_fifo/buff[0][6] , \i15/tx_fifo/buff[0][7] , \i15/tx_fifo/buff[1][0] , 
        \i15/tx_fifo/buff[1][1] , \i15/tx_fifo/buff[1][2] , \i15/tx_fifo/buff[1][3] , 
        \i15/tx_fifo/buff[1][4] , \i15/tx_fifo/buff[1][5] , \i15/tx_fifo/buff[1][6] , 
        \i15/tx_fifo/buff[1][7] , \i15/tx_fifo/buff[2][0] , \i15/tx_fifo/buff[2][1] , 
        \i15/tx_fifo/buff[2][2] , \i15/tx_fifo/buff[2][3] , \i15/tx_fifo/buff[2][4] , 
        \i15/tx_fifo/buff[2][5] , \i15/tx_fifo/buff[2][6] , \i15/tx_fifo/buff[2][7] , 
        \i15/tx_fifo/buff[3][0] , \i15/tx_fifo/buff[3][1] , \i15/tx_fifo/buff[3][2] , 
        \i15/tx_fifo/buff[3][3] , \i15/tx_fifo/buff[3][4] , \i15/tx_fifo/buff[3][5] , 
        \i15/tx_fifo/buff[3][6] , \i15/tx_fifo/buff[3][7] , \i15/tx_fifo/buff[4][0] , 
        \i15/tx_fifo/buff[4][1] , \i15/tx_fifo/buff[4][2] , \i15/tx_fifo/buff[4][3] , 
        \i15/tx_fifo/buff[4][4] , \i15/tx_fifo/buff[4][5] , \i15/tx_fifo/buff[4][6] , 
        \i15/tx_fifo/buff[4][7] , \i15/tx_fifo/buff[5][0] , \i15/tx_fifo/buff[5][1] , 
        \i15/tx_fifo/buff[5][2] , \i15/tx_fifo/buff[5][3] , \i15/tx_fifo/buff[5][4] , 
        \i15/tx_fifo/buff[5][5] , \i15/tx_fifo/buff[5][6] , \i15/tx_fifo/buff[5][7] , 
        \i15/tx_fifo/buff[6][0] , \i15/tx_fifo/buff[6][1] , \i15/tx_fifo/buff[6][2] , 
        \i15/tx_fifo/buff[6][3] , \i15/tx_fifo/buff[6][4] , \i15/tx_fifo/buff[6][5] , 
        \i15/tx_fifo/buff[6][6] , \i15/tx_fifo/buff[6][7] , \i15/tx_fifo/buff[7][0] , 
        \i15/tx_fifo/buff[7][1] , \i15/tx_fifo/buff[7][2] , \i15/tx_fifo/buff[7][3] , 
        \i15/tx_fifo/buff[7][4] , \i15/tx_fifo/buff[7][5] , \i15/tx_fifo/buff[7][6] , 
        \i15/tx_fifo/buff[7][7] , \i15/tx_fifo/buff[8][0] , \i15/tx_fifo/buff[8][1] , 
        \i15/tx_fifo/buff[8][2] , \i15/tx_fifo/buff[8][3] , \i15/tx_fifo/buff[8][4] , 
        \i15/tx_fifo/buff[8][5] , \i15/tx_fifo/buff[8][6] , \i15/tx_fifo/buff[8][7] , 
        \i15/tx_fifo/buff[9][0] , \i15/tx_fifo/buff[9][1] , \i15/tx_fifo/buff[9][2] , 
        \i15/tx_fifo/buff[9][3] , \i15/tx_fifo/buff[9][4] , \i15/tx_fifo/buff[9][5] , 
        \i15/tx_fifo/buff[9][6] , \i15/tx_fifo/buff[9][7] , \i15/tx_fifo/buff[10][0] , 
        \i15/tx_fifo/buff[10][1] , \i15/tx_fifo/buff[10][2] , \i15/tx_fifo/buff[10][3] , 
        \i15/tx_fifo/buff[10][4] , \i15/tx_fifo/buff[10][5] , \i15/tx_fifo/buff[10][6] , 
        \i15/tx_fifo/buff[10][7] , \i15/tx_fifo/buff[11][0] , \i15/tx_fifo/buff[11][1] , 
        \i15/tx_fifo/buff[11][2] , \i15/tx_fifo/buff[11][3] , \i15/tx_fifo/buff[11][4] , 
        \i15/tx_fifo/buff[11][5] , \i15/tx_fifo/buff[11][6] , \i15/tx_fifo/buff[11][7] , 
        \i15/tx_fifo/buff[12][0] , \i15/tx_fifo/buff[12][1] , \i15/tx_fifo/buff[12][2] , 
        \i15/tx_fifo/buff[12][3] , \i15/tx_fifo/buff[12][4] , \i15/tx_fifo/buff[12][5] , 
        \i15/tx_fifo/buff[12][6] , \i15/tx_fifo/buff[12][7] , \i15/tx_fifo/buff[13][0] , 
        \i15/tx_fifo/buff[13][1] , \i15/tx_fifo/buff[13][2] , \i15/tx_fifo/buff[13][3] , 
        \i15/tx_fifo/buff[13][4] , \i15/tx_fifo/buff[13][5] , \i15/tx_fifo/buff[13][6] , 
        \i15/tx_fifo/buff[13][7] , \i15/tx_fifo/buff[14][0] , \i15/tx_fifo/buff[14][1] , 
        \i15/tx_fifo/buff[14][2] , \i15/tx_fifo/buff[14][3] , \i15/tx_fifo/buff[14][4] , 
        \i15/tx_fifo/buff[14][5] , \i15/tx_fifo/buff[14][6] , \i15/tx_fifo/buff[14][7] , 
        \i15/tx_fifo/buff[15][0] , \i15/tx_fifo/buff[15][1] , \i15/tx_fifo/buff[15][2] , 
        \i15/tx_fifo/buff[15][3] , \i15/tx_fifo/buff[15][4] , \i15/tx_fifo/buff[15][5] , 
        \i15/tx_fifo/buff[15][6] , \i15/tx_fifo/buff[15][7] , \i15/tx_fifo/buff[16][0] , 
        \i15/tx_fifo/buff[16][1] , \i15/tx_fifo/buff[16][2] , \i15/tx_fifo/buff[16][3] , 
        \i15/tx_fifo/buff[16][4] , \i15/tx_fifo/buff[16][5] , \i15/tx_fifo/buff[16][6] , 
        \i15/tx_fifo/buff[16][7] , \i15/tx_fifo/buff[17][0] , \i15/tx_fifo/buff[17][1] , 
        \i15/tx_fifo/buff[17][2] , \i15/tx_fifo/buff[17][3] , \i15/tx_fifo/buff[17][4] , 
        \i15/tx_fifo/buff[17][5] , \i15/tx_fifo/buff[17][6] , \i15/tx_fifo/buff[17][7] , 
        \i15/tx_fifo/buff[18][0] , \i15/tx_fifo/buff[18][1] , \i15/tx_fifo/buff[18][2] , 
        \i15/tx_fifo/buff[18][3] , \i15/tx_fifo/buff[18][4] , \i15/tx_fifo/buff[18][5] , 
        \i15/tx_fifo/buff[18][6] , \i15/tx_fifo/buff[18][7] , \i15/tx_fifo/buff[19][0] , 
        \i15/tx_fifo/buff[19][1] , \i15/tx_fifo/buff[19][2] , \i15/tx_fifo/buff[19][3] , 
        \i15/tx_fifo/buff[19][4] , \i15/tx_fifo/buff[19][5] , \i15/tx_fifo/buff[19][6] , 
        \i15/tx_fifo/buff[19][7] , \i15/tx_fifo/buff[20][0] , \i15/tx_fifo/buff[20][1] , 
        \i15/tx_fifo/buff[20][2] , \i15/tx_fifo/buff[20][3] , \i15/tx_fifo/buff[20][4] , 
        \i15/tx_fifo/buff[20][5] , \i15/tx_fifo/buff[20][6] , \i15/tx_fifo/buff[20][7] , 
        \i15/tx_fifo/buff[21][0] , \i15/tx_fifo/buff[21][1] , \i15/tx_fifo/buff[21][2] , 
        \i15/tx_fifo/buff[21][3] , \i15/tx_fifo/buff[21][4] , \i15/tx_fifo/buff[21][5] , 
        \i15/tx_fifo/buff[21][6] , \i15/tx_fifo/buff[21][7] , \i15/tx_fifo/buff[22][0] , 
        \i15/tx_fifo/buff[22][1] , \i15/tx_fifo/buff[22][2] , \i15/tx_fifo/buff[22][3] , 
        \i15/tx_fifo/buff[22][4] , \i15/tx_fifo/buff[22][5] , \i15/tx_fifo/buff[22][6] , 
        \i15/tx_fifo/buff[22][7] , \i15/tx_fifo/buff[23][0] , \i15/tx_fifo/buff[23][1] , 
        \i15/tx_fifo/buff[23][2] , \i15/tx_fifo/buff[23][3] , \i15/tx_fifo/buff[23][4] , 
        \i15/tx_fifo/buff[23][5] , \i15/tx_fifo/buff[23][6] , \i15/tx_fifo/buff[23][7] , 
        \i15/tx_fifo/buff[24][0] , \i15/tx_fifo/buff[24][1] , \i15/tx_fifo/buff[24][2] , 
        \i15/tx_fifo/buff[24][3] , \i15/tx_fifo/buff[24][4] , \i15/tx_fifo/buff[24][5] , 
        \i15/tx_fifo/buff[24][6] , \i15/tx_fifo/buff[24][7] , \i15/tx_fifo/buff[25][0] , 
        \i15/tx_fifo/buff[25][1] , \i15/tx_fifo/buff[25][2] , \i15/tx_fifo/buff[25][3] , 
        \i15/tx_fifo/buff[25][4] , \i15/tx_fifo/buff[25][5] , \i15/tx_fifo/buff[25][6] , 
        \i15/tx_fifo/buff[25][7] , \i15/tx_fifo/buff[26][0] , \i15/tx_fifo/buff[26][1] , 
        \i15/tx_fifo/buff[26][2] , \i15/tx_fifo/buff[26][3] , \i15/tx_fifo/buff[26][4] , 
        \i15/tx_fifo/buff[26][5] , \i15/tx_fifo/buff[26][6] , \i15/tx_fifo/buff[26][7] , 
        \i15/tx_fifo/buff[27][0] , \i15/tx_fifo/buff[27][1] , \i15/tx_fifo/buff[27][2] , 
        \i15/tx_fifo/buff[27][3] , \i15/tx_fifo/buff[27][4] , \i15/tx_fifo/buff[27][5] , 
        \i15/tx_fifo/buff[27][6] , \i15/tx_fifo/buff[27][7] , \i15/tx_fifo/buff[28][0] , 
        \i15/tx_fifo/buff[28][1] , \i15/tx_fifo/buff[28][2] , \i15/tx_fifo/buff[28][3] , 
        \i15/tx_fifo/buff[28][4] , \i15/tx_fifo/buff[28][5] , \i15/tx_fifo/buff[28][6] , 
        \i15/tx_fifo/buff[28][7] , \i15/tx_fifo/buff[29][0] , \i15/tx_fifo/buff[29][1] , 
        \i15/tx_fifo/buff[29][2] , \i15/tx_fifo/buff[29][3] , \i15/tx_fifo/buff[29][4] , 
        \i15/tx_fifo/buff[29][5] , \i15/tx_fifo/buff[29][6] , \i15/tx_fifo/buff[29][7] , 
        \i15/tx_fifo/buff[30][0] , \i15/tx_fifo/buff[30][1] , \i15/tx_fifo/buff[30][2] , 
        \i15/tx_fifo/buff[30][3] , \i15/tx_fifo/buff[30][4] , \i15/tx_fifo/buff[30][5] , 
        \i15/tx_fifo/buff[30][6] , \i15/tx_fifo/buff[30][7] , \i15/tx_fifo/buff[31][0] , 
        \i15/tx_fifo/buff[31][1] , \i15/tx_fifo/buff[31][2] , \i15/tx_fifo/buff[31][3] , 
        \i15/tx_fifo/buff[31][4] , \i15/tx_fifo/buff[31][5] , \i15/tx_fifo/buff[31][6] , 
        \i15/tx_fifo/buff[31][7] , \i15/tx_fifo/buff[32][0] , \i15/tx_fifo/buff[32][1] , 
        \i15/tx_fifo/buff[32][2] , \i15/tx_fifo/buff[32][3] , \i15/tx_fifo/buff[32][4] , 
        \i15/tx_fifo/buff[32][5] , \i15/tx_fifo/buff[32][6] , \i15/tx_fifo/buff[32][7] , 
        \i15/tx_fifo/buff[33][0] , \i15/tx_fifo/buff[33][1] , \i15/tx_fifo/buff[33][2] , 
        \i15/tx_fifo/buff[33][3] , \i15/tx_fifo/buff[33][4] , \i15/tx_fifo/buff[33][5] , 
        \i15/tx_fifo/buff[33][6] , \i15/tx_fifo/buff[33][7] , \i15/tx_fifo/buff[34][0] , 
        \i15/tx_fifo/buff[34][1] , \i15/tx_fifo/buff[34][2] , \i15/tx_fifo/buff[34][3] , 
        \i15/tx_fifo/buff[34][4] , \i15/tx_fifo/buff[34][5] , \i15/tx_fifo/buff[34][6] , 
        \i15/tx_fifo/buff[34][7] , \i15/tx_fifo/buff[35][0] , \i15/tx_fifo/buff[35][1] , 
        \i15/tx_fifo/buff[35][2] , \i15/tx_fifo/buff[35][3] , \i15/tx_fifo/buff[35][4] , 
        \i15/tx_fifo/buff[35][5] , \i15/tx_fifo/buff[35][6] , \i15/tx_fifo/buff[35][7] , 
        \i15/tx_fifo/buff[36][0] , \i15/tx_fifo/buff[36][1] , \i15/tx_fifo/buff[36][2] , 
        \i15/tx_fifo/buff[36][3] , \i15/tx_fifo/buff[36][4] , \i15/tx_fifo/buff[36][5] , 
        \i15/tx_fifo/buff[36][6] , \i15/tx_fifo/buff[36][7] , \i15/tx_fifo/buff[37][0] , 
        \i15/tx_fifo/buff[37][1] , \i15/tx_fifo/buff[37][2] , \i15/tx_fifo/buff[37][3] , 
        \i15/tx_fifo/buff[37][4] , \i15/tx_fifo/buff[37][5] , \i15/tx_fifo/buff[37][6] , 
        \i15/tx_fifo/buff[37][7] , \i15/tx_fifo/buff[38][0] , \i15/tx_fifo/buff[38][1] , 
        \i15/tx_fifo/buff[38][2] , \i15/tx_fifo/buff[38][3] , \i15/tx_fifo/buff[38][4] , 
        \i15/tx_fifo/buff[38][5] , \i15/tx_fifo/buff[38][6] , \i15/tx_fifo/buff[38][7] , 
        \i15/tx_fifo/buff[39][0] , \i15/tx_fifo/buff[39][1] , \i15/tx_fifo/buff[39][2] , 
        \i15/tx_fifo/buff[39][3] , \i15/tx_fifo/buff[39][4] , \i15/tx_fifo/buff[39][5] , 
        \i15/tx_fifo/buff[39][6] , \i15/tx_fifo/buff[39][7] , \i15/tx_fifo/buff[40][0] , 
        \i15/tx_fifo/buff[40][1] , \i15/tx_fifo/buff[40][2] , \i15/tx_fifo/buff[40][3] , 
        \i15/tx_fifo/buff[40][4] , \i15/tx_fifo/buff[40][5] , \i15/tx_fifo/buff[40][6] , 
        \i15/tx_fifo/buff[40][7] , \i15/tx_fifo/buff[41][0] , \i15/tx_fifo/buff[41][1] , 
        \i15/tx_fifo/buff[41][2] , \i15/tx_fifo/buff[41][3] , \i15/tx_fifo/buff[41][4] , 
        \i15/tx_fifo/buff[41][5] , \i15/tx_fifo/buff[41][6] , \i15/tx_fifo/buff[41][7] , 
        \i15/tx_fifo/buff[42][0] , \i15/tx_fifo/buff[42][1] , \i15/tx_fifo/buff[42][2] , 
        \i15/tx_fifo/buff[42][3] , \i15/tx_fifo/buff[42][4] , \i15/tx_fifo/buff[42][5] , 
        \i15/tx_fifo/buff[42][6] , \i15/tx_fifo/buff[42][7] , \i15/tx_fifo/buff[43][0] , 
        \i15/tx_fifo/buff[43][1] , \i15/tx_fifo/buff[43][2] , \i15/tx_fifo/buff[43][3] , 
        \i15/tx_fifo/buff[43][4] , \i15/tx_fifo/buff[43][5] , \i15/tx_fifo/buff[43][6] , 
        \i15/tx_fifo/buff[43][7] , \i15/tx_fifo/buff[44][0] , \i15/tx_fifo/buff[44][1] , 
        \i15/tx_fifo/buff[44][2] , \i15/tx_fifo/buff[44][3] , \i15/tx_fifo/buff[44][4] , 
        \i15/tx_fifo/buff[44][5] , \i15/tx_fifo/buff[44][6] , \i15/tx_fifo/buff[44][7] , 
        \i15/tx_fifo/buff[45][0] , \i15/tx_fifo/buff[45][1] , \i15/tx_fifo/buff[45][2] , 
        \i15/tx_fifo/buff[45][3] , \i15/tx_fifo/buff[45][4] , \i15/tx_fifo/buff[45][5] , 
        \i15/tx_fifo/buff[45][6] , \i15/tx_fifo/buff[45][7] , \i15/tx_fifo/buff[46][0] , 
        \i15/tx_fifo/buff[46][1] , \i15/tx_fifo/buff[46][2] , \i15/tx_fifo/buff[46][3] , 
        \i15/tx_fifo/buff[46][4] , \i15/tx_fifo/buff[46][5] , \i15/tx_fifo/buff[46][6] , 
        \i15/tx_fifo/buff[46][7] , \i15/tx_fifo/buff[47][0] , \i15/tx_fifo/buff[47][1] , 
        \i15/tx_fifo/buff[47][2] , \i15/tx_fifo/buff[47][3] , \i15/tx_fifo/buff[47][4] , 
        \i15/tx_fifo/buff[47][5] , \i15/tx_fifo/buff[47][6] , \i15/tx_fifo/buff[47][7] , 
        \i15/tx_fifo/buff[48][0] , \i15/tx_fifo/buff[48][1] , \i15/tx_fifo/buff[48][2] , 
        \i15/tx_fifo/buff[48][3] , \i15/tx_fifo/buff[48][4] , \i15/tx_fifo/buff[48][5] , 
        \i15/tx_fifo/buff[48][6] , \i15/tx_fifo/buff[48][7] , \i15/tx_fifo/buff[49][0] , 
        \i15/tx_fifo/buff[49][1] , \i15/tx_fifo/buff[49][2] , \i15/tx_fifo/buff[49][3] , 
        \i15/tx_fifo/buff[49][4] , \i15/tx_fifo/buff[49][5] , \i15/tx_fifo/buff[49][6] , 
        \i15/tx_fifo/buff[49][7] , \i15/tx_fifo/buff[50][0] , \i15/tx_fifo/buff[50][1] , 
        \i15/tx_fifo/buff[50][2] , \i15/tx_fifo/buff[50][3] , \i15/tx_fifo/buff[50][4] , 
        \i15/tx_fifo/buff[50][5] , \i15/tx_fifo/buff[50][6] , \i15/tx_fifo/buff[50][7] , 
        \i15/tx_fifo/buff[51][0] , \i15/tx_fifo/buff[51][1] , \i15/tx_fifo/buff[51][2] , 
        \i15/tx_fifo/buff[51][3] , \i15/tx_fifo/buff[51][4] , \i15/tx_fifo/buff[51][5] , 
        \i15/tx_fifo/buff[51][6] , \i15/tx_fifo/buff[51][7] , \i15/tx_fifo/buff[52][0] , 
        \i15/tx_fifo/buff[52][1] , \i15/tx_fifo/buff[52][2] , \i15/tx_fifo/buff[52][3] , 
        \i15/tx_fifo/buff[52][4] , \i15/tx_fifo/buff[52][5] , \i15/tx_fifo/buff[52][6] , 
        \i15/tx_fifo/buff[52][7] , \i15/tx_fifo/buff[53][0] , \i15/tx_fifo/buff[53][1] , 
        \i15/tx_fifo/buff[53][2] , \i15/tx_fifo/buff[53][3] , \i15/tx_fifo/buff[53][4] , 
        \i15/tx_fifo/buff[53][5] , \i15/tx_fifo/buff[53][6] , \i15/tx_fifo/buff[53][7] , 
        \i15/tx_fifo/buff[54][0] , \i15/tx_fifo/buff[54][1] , \i15/tx_fifo/buff[54][2] , 
        \i15/tx_fifo/buff[54][3] , \i15/tx_fifo/buff[54][4] , \i15/tx_fifo/buff[54][5] , 
        \i15/tx_fifo/buff[54][6] , \i15/tx_fifo/buff[54][7] , \i15/tx_fifo/buff[55][0] , 
        \i15/tx_fifo/buff[55][1] , \i15/tx_fifo/buff[55][2] , \i15/tx_fifo/buff[55][3] , 
        \i15/tx_fifo/buff[55][4] , \i15/tx_fifo/buff[55][5] , \i15/tx_fifo/buff[55][6] , 
        \i15/tx_fifo/buff[55][7] , \i15/tx_fifo/buff[56][0] , \i15/tx_fifo/buff[56][1] , 
        \i15/tx_fifo/buff[56][2] , \i15/tx_fifo/buff[56][3] , \i15/tx_fifo/buff[56][4] , 
        \i15/tx_fifo/buff[56][5] , \i15/tx_fifo/buff[56][6] , \i15/tx_fifo/buff[56][7] , 
        \i15/tx_fifo/buff[57][0] , \i15/tx_fifo/buff[57][1] , \i15/tx_fifo/buff[57][2] , 
        \i15/tx_fifo/buff[57][3] , \i15/tx_fifo/buff[57][4] , \i15/tx_fifo/buff[57][5] , 
        \i15/tx_fifo/buff[57][6] , \i15/tx_fifo/buff[57][7] , \i15/tx_fifo/buff[58][0] , 
        \i15/tx_fifo/buff[58][1] , \i15/tx_fifo/buff[58][2] , \i15/tx_fifo/buff[58][3] , 
        \i15/tx_fifo/buff[58][4] , \i15/tx_fifo/buff[58][5] , \i15/tx_fifo/buff[58][6] , 
        \i15/tx_fifo/buff[58][7] , \i15/tx_fifo/buff[59][0] , \i15/tx_fifo/buff[59][1] , 
        \i15/tx_fifo/buff[59][2] , \i15/tx_fifo/buff[59][3] , \i15/tx_fifo/buff[59][4] , 
        \i15/tx_fifo/buff[59][5] , \i15/tx_fifo/buff[59][6] , \i15/tx_fifo/buff[59][7] , 
        \i15/tx_fifo/buff[60][0] , \i15/tx_fifo/buff[60][1] , \i15/tx_fifo/buff[60][2] , 
        \i15/tx_fifo/buff[60][3] , \i15/tx_fifo/buff[60][4] , \i15/tx_fifo/buff[60][5] , 
        \i15/tx_fifo/buff[60][6] , \i15/tx_fifo/buff[60][7] , \i15/tx_fifo/buff[61][0] , 
        \i15/tx_fifo/buff[61][1] , \i15/tx_fifo/buff[61][2] , \i15/tx_fifo/buff[61][3] , 
        \i15/tx_fifo/buff[61][4] , \i15/tx_fifo/buff[61][5] , \i15/tx_fifo/buff[61][6] , 
        \i15/tx_fifo/buff[61][7] , \i15/tx_fifo/buff[62][0] , \i15/tx_fifo/buff[62][1] , 
        \i15/tx_fifo/buff[62][2] , \i15/tx_fifo/buff[62][3] , \i15/tx_fifo/buff[62][4] , 
        \i15/tx_fifo/buff[62][5] , \i15/tx_fifo/buff[62][6] , \i15/tx_fifo/buff[62][7] , 
        \i15/tx_fifo/buff[63][0] , \i15/tx_fifo/buff[63][1] , \i15/tx_fifo/buff[63][2] , 
        \i15/tx_fifo/buff[63][3] , \i15/tx_fifo/buff[63][4] , \i15/tx_fifo/buff[63][5] , 
        \i15/tx_fifo/buff[63][6] , \i15/tx_fifo/buff[63][7] , \i15/tx_fifo/buff[64][0] , 
        \i15/tx_fifo/buff[64][1] , \i15/tx_fifo/buff[64][2] , \i15/tx_fifo/buff[64][3] , 
        \i15/tx_fifo/buff[64][4] , \i15/tx_fifo/buff[64][5] , \i15/tx_fifo/buff[64][6] , 
        \i15/tx_fifo/buff[64][7] , \i15/tx_fifo/buff[65][0] , \i15/tx_fifo/buff[65][1] , 
        \i15/tx_fifo/buff[65][2] , \i15/tx_fifo/buff[65][3] , \i15/tx_fifo/buff[65][4] , 
        \i15/tx_fifo/buff[65][5] , \i15/tx_fifo/buff[65][6] , \i15/tx_fifo/buff[65][7] , 
        \i15/tx_fifo/buff[66][0] , \i15/tx_fifo/buff[66][1] , \i15/tx_fifo/buff[66][2] , 
        \i15/tx_fifo/buff[66][3] , \i15/tx_fifo/buff[66][4] , \i15/tx_fifo/buff[66][5] , 
        \i15/tx_fifo/buff[66][6] , \i15/tx_fifo/buff[66][7] , \i15/tx_fifo/buff[67][0] , 
        \i15/tx_fifo/buff[67][1] , \i15/tx_fifo/buff[67][2] , \i15/tx_fifo/buff[67][3] , 
        \i15/tx_fifo/buff[67][4] , \i15/tx_fifo/buff[67][5] , \i15/tx_fifo/buff[67][6] , 
        \i15/tx_fifo/buff[67][7] , \i15/tx_fifo/buff[68][0] , \i15/tx_fifo/buff[68][1] , 
        \i15/tx_fifo/buff[68][2] , \i15/tx_fifo/buff[68][3] , \i15/tx_fifo/buff[68][4] , 
        \i15/tx_fifo/buff[68][5] , \i15/tx_fifo/buff[68][6] , \i15/tx_fifo/buff[68][7] , 
        \i15/tx_fifo/buff[69][0] , \i15/tx_fifo/buff[69][1] , \i15/tx_fifo/buff[69][2] , 
        \i15/tx_fifo/buff[69][3] , \i15/tx_fifo/buff[69][4] , \i15/tx_fifo/buff[69][5] , 
        \i15/tx_fifo/buff[69][6] , \i15/tx_fifo/buff[69][7] , \i15/tx_fifo/buff[70][0] , 
        \i15/tx_fifo/buff[70][1] , \i15/tx_fifo/buff[70][2] , \i15/tx_fifo/buff[70][3] , 
        \i15/tx_fifo/buff[70][4] , \i15/tx_fifo/buff[70][5] , \i15/tx_fifo/buff[70][6] , 
        \i15/tx_fifo/buff[70][7] , \i15/tx_fifo/buff[71][0] , \i15/tx_fifo/buff[71][1] , 
        \i15/tx_fifo/buff[71][2] , \i15/tx_fifo/buff[71][3] , \i15/tx_fifo/buff[71][4] , 
        \i15/tx_fifo/buff[71][5] , \i15/tx_fifo/buff[71][6] , \i15/tx_fifo/buff[71][7] , 
        \i15/tx_fifo/buff[72][0] , \i15/tx_fifo/buff[72][1] , \i15/tx_fifo/buff[72][2] , 
        \i15/tx_fifo/buff[72][3] , \i15/tx_fifo/buff[72][4] , \i15/tx_fifo/buff[72][5] , 
        \i15/tx_fifo/buff[72][6] , \i15/tx_fifo/buff[72][7] , \i15/tx_fifo/buff[73][0] , 
        \i15/tx_fifo/buff[73][1] , \i15/tx_fifo/buff[73][2] , \i15/tx_fifo/buff[73][3] , 
        \i15/tx_fifo/buff[73][4] , \i15/tx_fifo/buff[73][5] , \i15/tx_fifo/buff[73][6] , 
        \i15/tx_fifo/buff[73][7] , \i15/tx_fifo/buff[74][0] , \i15/tx_fifo/buff[74][1] , 
        \i15/tx_fifo/buff[74][2] , \i15/tx_fifo/buff[74][3] , \i15/tx_fifo/buff[74][4] , 
        \i15/tx_fifo/buff[74][5] , \i15/tx_fifo/buff[74][6] , \i15/tx_fifo/buff[74][7] , 
        \i15/tx_fifo/buff[75][0] , \i15/tx_fifo/buff[75][1] , \i15/tx_fifo/buff[75][2] , 
        \i15/tx_fifo/buff[75][3] , \i15/tx_fifo/buff[75][4] , \i15/tx_fifo/buff[75][5] , 
        \i15/tx_fifo/buff[75][6] , \i15/tx_fifo/buff[75][7] , \i15/tx_fifo/buff[76][0] , 
        \i15/tx_fifo/buff[76][1] , \i15/tx_fifo/buff[76][2] , \i15/tx_fifo/buff[76][3] , 
        \i15/tx_fifo/buff[76][4] , \i15/tx_fifo/buff[76][5] , \i15/tx_fifo/buff[76][6] , 
        \i15/tx_fifo/buff[76][7] , \i15/tx_fifo/buff[77][0] , \i15/tx_fifo/buff[77][1] , 
        \i15/tx_fifo/buff[77][2] , \i15/tx_fifo/buff[77][3] , \i15/tx_fifo/buff[77][4] , 
        \i15/tx_fifo/buff[77][5] , \i15/tx_fifo/buff[77][6] , \i15/tx_fifo/buff[77][7] , 
        \i15/tx_fifo/buff[78][0] , \i15/tx_fifo/buff[78][1] , \i15/tx_fifo/buff[78][2] , 
        \i15/tx_fifo/buff[78][3] , \i15/tx_fifo/buff[78][4] , \i15/tx_fifo/buff[78][5] , 
        \i15/tx_fifo/buff[78][6] , \i15/tx_fifo/buff[78][7] , \i15/tx_fifo/buff[79][0] , 
        \i15/tx_fifo/buff[79][1] , \i15/tx_fifo/buff[79][2] , \i15/tx_fifo/buff[79][3] , 
        \i15/tx_fifo/buff[79][4] , \i15/tx_fifo/buff[79][5] , \i15/tx_fifo/buff[79][6] , 
        \i15/tx_fifo/buff[79][7] , \i15/tx_fifo/buff[80][0] , \i15/tx_fifo/buff[80][1] , 
        \i15/tx_fifo/buff[80][2] , \i15/tx_fifo/buff[80][3] , \i15/tx_fifo/buff[80][4] , 
        \i15/tx_fifo/buff[80][5] , \i15/tx_fifo/buff[80][6] , \i15/tx_fifo/buff[80][7] , 
        \i15/tx_fifo/buff[81][0] , \i15/tx_fifo/buff[81][1] , \i15/tx_fifo/buff[81][2] , 
        \i15/tx_fifo/buff[81][3] , \i15/tx_fifo/buff[81][4] , \i15/tx_fifo/buff[81][5] , 
        \i15/tx_fifo/buff[81][6] , \i15/tx_fifo/buff[81][7] , \i15/tx_fifo/buff[82][0] , 
        \i15/tx_fifo/buff[82][1] , \i15/tx_fifo/buff[82][2] , \i15/tx_fifo/buff[82][3] , 
        \i15/tx_fifo/buff[82][4] , \i15/tx_fifo/buff[82][5] , \i15/tx_fifo/buff[82][6] , 
        \i15/tx_fifo/buff[82][7] , \i15/tx_fifo/buff[83][0] , \i15/tx_fifo/buff[83][1] , 
        \i15/tx_fifo/buff[83][2] , \i15/tx_fifo/buff[83][3] , \i15/tx_fifo/buff[83][4] , 
        \i15/tx_fifo/buff[83][5] , \i15/tx_fifo/buff[83][6] , \i15/tx_fifo/buff[83][7] , 
        \i15/tx_fifo/buff[84][0] , \i15/tx_fifo/buff[84][1] , \i15/tx_fifo/buff[84][2] , 
        \i15/tx_fifo/buff[84][3] , \i15/tx_fifo/buff[84][4] , \i15/tx_fifo/buff[84][5] , 
        \i15/tx_fifo/buff[84][6] , \i15/tx_fifo/buff[84][7] , \i15/tx_fifo/buff[85][0] , 
        \i15/tx_fifo/buff[85][1] , \i15/tx_fifo/buff[85][2] , \i15/tx_fifo/buff[85][3] , 
        \i15/tx_fifo/buff[85][4] , \i15/tx_fifo/buff[85][5] , \i15/tx_fifo/buff[85][6] , 
        \i15/tx_fifo/buff[85][7] , \i15/tx_fifo/buff[86][0] , \i15/tx_fifo/buff[86][1] , 
        \i15/tx_fifo/buff[86][2] , \i15/tx_fifo/buff[86][3] , \i15/tx_fifo/buff[86][4] , 
        \i15/tx_fifo/buff[86][5] , \i15/tx_fifo/buff[86][6] , \i15/tx_fifo/buff[86][7] , 
        \i15/tx_fifo/buff[87][0] , \i15/tx_fifo/buff[87][1] , \i15/tx_fifo/buff[87][2] , 
        \i15/tx_fifo/buff[87][3] , \i15/tx_fifo/buff[87][4] , \i15/tx_fifo/buff[87][5] , 
        \i15/tx_fifo/buff[87][6] , \i15/tx_fifo/buff[87][7] , \i15/tx_fifo/buff[88][0] , 
        \i15/tx_fifo/buff[88][1] , \i15/tx_fifo/buff[88][2] , \i15/tx_fifo/buff[88][3] , 
        \i15/tx_fifo/buff[88][4] , \i15/tx_fifo/buff[88][5] , \i15/tx_fifo/buff[88][6] , 
        \i15/tx_fifo/buff[88][7] , \i15/tx_fifo/buff[89][0] , \i15/tx_fifo/buff[89][1] , 
        \i15/tx_fifo/buff[89][2] , \i15/tx_fifo/buff[89][3] , \i15/tx_fifo/buff[89][4] , 
        \i15/tx_fifo/buff[89][5] , \i15/tx_fifo/buff[89][6] , \i15/tx_fifo/buff[89][7] , 
        \i15/tx_fifo/buff[90][0] , \i15/tx_fifo/buff[90][1] , \i15/tx_fifo/buff[90][2] , 
        \i15/tx_fifo/buff[90][3] , \i15/tx_fifo/buff[90][4] , \i15/tx_fifo/buff[90][5] , 
        \i15/tx_fifo/buff[90][6] , \i15/tx_fifo/buff[90][7] , \i15/tx_fifo/buff[91][0] , 
        \i15/tx_fifo/buff[91][1] , \i15/tx_fifo/buff[91][2] , \i15/tx_fifo/buff[91][3] , 
        \i15/tx_fifo/buff[91][4] , \i15/tx_fifo/buff[91][5] , \i15/tx_fifo/buff[91][6] , 
        \i15/tx_fifo/buff[91][7] , \i15/tx_fifo/buff[92][0] , \i15/tx_fifo/buff[92][1] , 
        \i15/tx_fifo/buff[92][2] , \i15/tx_fifo/buff[92][3] , \i15/tx_fifo/buff[92][4] , 
        \i15/tx_fifo/buff[92][5] , \i15/tx_fifo/buff[92][6] , \i15/tx_fifo/buff[92][7] , 
        \i15/tx_fifo/buff[93][0] , \i15/tx_fifo/buff[93][1] , \i15/tx_fifo/buff[93][2] , 
        \i15/tx_fifo/buff[93][3] , \i15/tx_fifo/buff[93][4] , \i15/tx_fifo/buff[93][5] , 
        \i15/tx_fifo/buff[93][6] , \i15/tx_fifo/buff[93][7] , \i15/tx_fifo/buff[94][0] , 
        \i15/tx_fifo/buff[94][1] , \i15/tx_fifo/buff[94][2] , \i15/tx_fifo/buff[94][3] , 
        \i15/tx_fifo/buff[94][4] , \i15/tx_fifo/buff[94][5] , \i15/tx_fifo/buff[94][6] , 
        \i15/tx_fifo/buff[94][7] , \i15/tx_fifo/buff[95][0] , \i15/tx_fifo/buff[95][1] , 
        \i15/tx_fifo/buff[95][2] , \i15/tx_fifo/buff[95][3] , \i15/tx_fifo/buff[95][4] , 
        \i15/tx_fifo/buff[95][5] , \i15/tx_fifo/buff[95][6] , \i15/tx_fifo/buff[95][7] , 
        \i15/tx_fifo/buff[96][0] , \i15/tx_fifo/buff[96][1] , \i15/tx_fifo/buff[96][2] , 
        \i15/tx_fifo/buff[96][3] , \i15/tx_fifo/buff[96][4] , \i15/tx_fifo/buff[96][5] , 
        \i15/tx_fifo/buff[96][6] , \i15/tx_fifo/buff[96][7] , \i15/tx_fifo/buff[97][0] , 
        \i15/tx_fifo/buff[97][1] , \i15/tx_fifo/buff[97][2] , \i15/tx_fifo/buff[97][3] , 
        \i15/tx_fifo/buff[97][4] , \i15/tx_fifo/buff[97][5] , \i15/tx_fifo/buff[97][6] , 
        \i15/tx_fifo/buff[97][7] , \i15/tx_fifo/buff[98][0] , \i15/tx_fifo/buff[98][1] , 
        \i15/tx_fifo/buff[98][2] , \i15/tx_fifo/buff[98][3] , \i15/tx_fifo/buff[98][4] , 
        \i15/tx_fifo/buff[98][5] , \i15/tx_fifo/buff[98][6] , \i15/tx_fifo/buff[98][7] , 
        \i15/tx_fifo/buff[99][0] , \i15/tx_fifo/buff[99][1] , \i15/tx_fifo/buff[99][2] , 
        \i15/tx_fifo/buff[99][3] , \i15/tx_fifo/buff[99][4] , \i15/tx_fifo/buff[99][5] , 
        \i15/tx_fifo/buff[99][6] , \i15/tx_fifo/buff[99][7] , \i15/tx_fifo/buff[100][0] , 
        \i15/tx_fifo/buff[100][1] , \i15/tx_fifo/buff[100][2] , \i15/tx_fifo/buff[100][3] , 
        \i15/tx_fifo/buff[100][4] , \i15/tx_fifo/buff[100][5] , \i15/tx_fifo/buff[100][6] , 
        \i15/tx_fifo/buff[100][7] , \i15/tx_fifo/buff[101][0] , \i15/tx_fifo/buff[101][1] , 
        \i15/tx_fifo/buff[101][2] , \i15/tx_fifo/buff[101][3] , \i15/tx_fifo/buff[101][4] , 
        \i15/tx_fifo/buff[101][5] , \i15/tx_fifo/buff[101][6] , \i15/tx_fifo/buff[101][7] , 
        \i15/tx_fifo/buff[102][0] , \i15/tx_fifo/buff[102][1] , \i15/tx_fifo/buff[102][2] , 
        \i15/tx_fifo/buff[102][3] , \i15/tx_fifo/buff[102][4] , \i15/tx_fifo/buff[102][5] , 
        \i15/tx_fifo/buff[102][6] , \i15/tx_fifo/buff[102][7] , \i15/tx_fifo/buff[103][0] , 
        \i15/tx_fifo/buff[103][1] , \i15/tx_fifo/buff[103][2] , \i15/tx_fifo/buff[103][3] , 
        \i15/tx_fifo/buff[103][4] , \i15/tx_fifo/buff[103][5] , \i15/tx_fifo/buff[103][6] , 
        \i15/tx_fifo/buff[103][7] , \i15/tx_fifo/buff[104][0] , \i15/tx_fifo/buff[104][1] , 
        \i15/tx_fifo/buff[104][2] , \i15/tx_fifo/buff[104][3] , \i15/tx_fifo/buff[104][4] , 
        \i15/tx_fifo/buff[104][5] , \i15/tx_fifo/buff[104][6] , \i15/tx_fifo/buff[104][7] , 
        \i15/tx_fifo/buff[105][0] , \i15/tx_fifo/buff[105][1] , \i15/tx_fifo/buff[105][2] , 
        \i15/tx_fifo/buff[105][3] , \i15/tx_fifo/buff[105][4] , \i15/tx_fifo/buff[105][5] , 
        \i15/tx_fifo/buff[105][6] , \i15/tx_fifo/buff[105][7] , \i15/tx_fifo/buff[106][0] , 
        \i15/tx_fifo/buff[106][1] , \i15/tx_fifo/buff[106][2] , \i15/tx_fifo/buff[106][3] , 
        \i15/tx_fifo/buff[106][4] , \i15/tx_fifo/buff[106][5] , \i15/tx_fifo/buff[106][6] , 
        \i15/tx_fifo/buff[106][7] , \i15/tx_fifo/buff[107][0] , \i15/tx_fifo/buff[107][1] , 
        \i15/tx_fifo/buff[107][2] , \i15/tx_fifo/buff[107][3] , \i15/tx_fifo/buff[107][4] , 
        \i15/tx_fifo/buff[107][5] , \i15/tx_fifo/buff[107][6] , \i15/tx_fifo/buff[107][7] , 
        \i15/tx_fifo/buff[108][0] , \i15/tx_fifo/buff[108][1] , \i15/tx_fifo/buff[108][2] , 
        \i15/tx_fifo/buff[108][3] , \i15/tx_fifo/buff[108][4] , \i15/tx_fifo/buff[108][5] , 
        \i15/tx_fifo/buff[108][6] , \i15/tx_fifo/buff[108][7] , \i15/tx_fifo/buff[109][0] , 
        \i15/tx_fifo/buff[109][1] , \i15/tx_fifo/buff[109][2] , \i15/tx_fifo/buff[109][3] , 
        \i15/tx_fifo/buff[109][4] , \i15/tx_fifo/buff[109][5] , \i15/tx_fifo/buff[109][6] , 
        \i15/tx_fifo/buff[109][7] , \i15/tx_fifo/buff[110][0] , \i15/tx_fifo/buff[110][1] , 
        \i15/tx_fifo/buff[110][2] , \i15/tx_fifo/buff[110][3] , \i15/tx_fifo/buff[110][4] , 
        \i15/tx_fifo/buff[110][5] , \i15/tx_fifo/buff[110][6] , \i15/tx_fifo/buff[110][7] , 
        \i15/tx_fifo/buff[111][0] , \i15/tx_fifo/buff[111][1] , \i15/tx_fifo/buff[111][2] , 
        \i15/tx_fifo/buff[111][3] , \i15/tx_fifo/buff[111][4] , \i15/tx_fifo/buff[111][5] , 
        \i15/tx_fifo/buff[111][6] , \i15/tx_fifo/buff[111][7] , \i15/tx_fifo/buff[112][0] , 
        \i15/tx_fifo/buff[112][1] , \i15/tx_fifo/buff[112][2] , \i15/tx_fifo/buff[112][3] , 
        \i15/tx_fifo/buff[112][4] , \i15/tx_fifo/buff[112][5] , \i15/tx_fifo/buff[112][6] , 
        \i15/tx_fifo/buff[112][7] , \i15/tx_fifo/buff[113][0] , \i15/tx_fifo/buff[113][1] , 
        \i15/tx_fifo/buff[113][2] , \i15/tx_fifo/buff[113][3] , \i15/tx_fifo/buff[113][4] , 
        \i15/tx_fifo/buff[113][5] , \i15/tx_fifo/buff[113][6] , \i15/tx_fifo/buff[113][7] , 
        \i15/tx_fifo/buff[114][0] , \i15/tx_fifo/buff[114][1] , \i15/tx_fifo/buff[114][2] , 
        \i15/tx_fifo/buff[114][3] , \i15/tx_fifo/buff[114][4] , \i15/tx_fifo/buff[114][5] , 
        \i15/tx_fifo/buff[114][6] , \i15/tx_fifo/buff[114][7] , \i15/tx_fifo/buff[115][0] , 
        \i15/tx_fifo/buff[115][1] , \i15/tx_fifo/buff[115][2] , \i15/tx_fifo/buff[115][3] , 
        \i15/tx_fifo/buff[115][4] , \i15/tx_fifo/buff[115][5] , \i15/tx_fifo/buff[115][6] , 
        \i15/tx_fifo/buff[115][7] , \i15/tx_fifo/buff[116][0] , \i15/tx_fifo/buff[116][1] , 
        \i15/tx_fifo/buff[116][2] , \i15/tx_fifo/buff[116][3] , \i15/tx_fifo/buff[116][4] , 
        \i15/tx_fifo/buff[116][5] , \i15/tx_fifo/buff[116][6] , \i15/tx_fifo/buff[116][7] , 
        \i15/tx_fifo/buff[117][0] , \i15/tx_fifo/buff[117][1] , \i15/tx_fifo/buff[117][2] , 
        \i15/tx_fifo/buff[117][3] , \i15/tx_fifo/buff[117][4] , \i15/tx_fifo/buff[117][5] , 
        \i15/tx_fifo/buff[117][6] , \i15/tx_fifo/buff[117][7] , \i15/tx_fifo/buff[118][0] , 
        \i15/tx_fifo/buff[118][1] , \i15/tx_fifo/buff[118][2] , \i15/tx_fifo/buff[118][3] , 
        \i15/tx_fifo/buff[118][4] , \i15/tx_fifo/buff[118][5] , \i15/tx_fifo/buff[118][6] , 
        \i15/tx_fifo/buff[118][7] , \i15/tx_fifo/buff[119][0] , \i15/tx_fifo/buff[119][1] , 
        \i15/tx_fifo/buff[119][2] , \i15/tx_fifo/buff[119][3] , \i15/tx_fifo/buff[119][4] , 
        \i15/tx_fifo/buff[119][5] , \i15/tx_fifo/buff[119][6] , \i15/tx_fifo/buff[119][7] , 
        \i15/tx_fifo/buff[120][0] , \i15/tx_fifo/buff[120][1] , \i15/tx_fifo/buff[120][2] , 
        \i15/tx_fifo/buff[120][3] , \i15/tx_fifo/buff[120][4] , \i15/tx_fifo/buff[120][5] , 
        \i15/tx_fifo/buff[120][6] , \i15/tx_fifo/buff[120][7] , \i15/tx_fifo/buff[121][0] , 
        \i15/tx_fifo/buff[121][1] , \i15/tx_fifo/buff[121][2] , \i15/tx_fifo/buff[121][3] , 
        \i15/tx_fifo/buff[121][4] , \i15/tx_fifo/buff[121][5] , \i15/tx_fifo/buff[121][6] , 
        \i15/tx_fifo/buff[121][7] , \i15/tx_fifo/buff[122][0] , \i15/tx_fifo/buff[122][1] , 
        \i15/tx_fifo/buff[122][2] , \i15/tx_fifo/buff[122][3] , \i15/tx_fifo/buff[122][4] , 
        \i15/tx_fifo/buff[122][5] , \i15/tx_fifo/buff[122][6] , \i15/tx_fifo/buff[122][7] , 
        \i15/tx_fifo/buff[123][0] , \i15/tx_fifo/buff[123][1] , \i15/tx_fifo/buff[123][2] , 
        \i15/tx_fifo/buff[123][3] , \i15/tx_fifo/buff[123][4] , \i15/tx_fifo/buff[123][5] , 
        \i15/tx_fifo/buff[123][6] , \i15/tx_fifo/buff[123][7] , \i15/tx_fifo/buff[124][0] , 
        \i15/tx_fifo/buff[124][1] , \i15/tx_fifo/buff[124][2] , \i15/tx_fifo/buff[124][3] , 
        \i15/tx_fifo/buff[124][4] , \i15/tx_fifo/buff[124][5] , \i15/tx_fifo/buff[124][6] , 
        \i15/tx_fifo/buff[124][7] , \i15/tx_fifo/buff[125][0] , \i15/tx_fifo/buff[125][1] , 
        \i15/tx_fifo/buff[125][2] , \i15/tx_fifo/buff[125][3] , \i15/tx_fifo/buff[125][4] , 
        \i15/tx_fifo/buff[125][5] , \i15/tx_fifo/buff[125][6] , \i15/tx_fifo/buff[125][7] , 
        \i15/tx_fifo/buff[126][0] , \i15/tx_fifo/buff[126][1] , \i15/tx_fifo/buff[126][2] , 
        \i15/tx_fifo/buff[126][3] , \i15/tx_fifo/buff[126][4] , \i15/tx_fifo/buff[126][5] , 
        \i15/tx_fifo/buff[126][6] , \i15/tx_fifo/buff[126][7] , \i15/tx_fifo/buff[127][0] , 
        \i15/tx_fifo/buff[127][1] , \i15/tx_fifo/buff[127][2] , \i15/tx_fifo/buff[127][3] , 
        \i15/tx_fifo/buff[127][4] , \i15/tx_fifo/buff[127][5] , \i15/tx_fifo/buff[127][6] , 
        \i15/tx_fifo/buff[127][7] , \i16/rx_fifo/buff[0][0] , \i16/rx_fifo/buff[0][1] , 
        \i16/rx_fifo/buff[0][2] , \i16/rx_fifo/buff[0][3] , \i16/rx_fifo/buff[0][4] , 
        \i16/rx_fifo/buff[0][5] , \i16/rx_fifo/buff[0][6] , \i16/rx_fifo/buff[0][7] , 
        \i16/rx_fifo/buff[1][0] , \i16/rx_fifo/buff[1][1] , \i16/rx_fifo/buff[1][2] , 
        \i16/rx_fifo/buff[1][3] , \i16/rx_fifo/buff[1][4] , \i16/rx_fifo/buff[1][5] , 
        \i16/rx_fifo/buff[1][6] , \i16/rx_fifo/buff[1][7] , \i16/rx_fifo/buff[2][0] , 
        \i16/rx_fifo/buff[2][1] , \i16/rx_fifo/buff[2][2] , \i16/rx_fifo/buff[2][3] , 
        \i16/rx_fifo/buff[2][4] , \i16/rx_fifo/buff[2][5] , \i16/rx_fifo/buff[2][6] , 
        \i16/rx_fifo/buff[2][7] , \i16/rx_fifo/buff[3][0] , \i16/rx_fifo/buff[3][1] , 
        \i16/rx_fifo/buff[3][2] , \i16/rx_fifo/buff[3][3] , \i16/rx_fifo/buff[3][4] , 
        \i16/rx_fifo/buff[3][5] , \i16/rx_fifo/buff[3][6] , \i16/rx_fifo/buff[3][7] , 
        \i16/rx_fifo/buff[4][0] , \i16/rx_fifo/buff[4][1] , \i16/rx_fifo/buff[4][2] , 
        \i16/rx_fifo/buff[4][3] , \i16/rx_fifo/buff[4][4] , \i16/rx_fifo/buff[4][5] , 
        \i16/rx_fifo/buff[4][6] , \i16/rx_fifo/buff[4][7] , \i16/rx_fifo/buff[5][0] , 
        \i16/rx_fifo/buff[5][1] , \i16/rx_fifo/buff[5][2] , \i16/rx_fifo/buff[5][3] , 
        \i16/rx_fifo/buff[5][4] , \i16/rx_fifo/buff[5][5] , \i16/rx_fifo/buff[5][6] , 
        \i16/rx_fifo/buff[5][7] , \i16/rx_fifo/buff[6][0] , \i16/rx_fifo/buff[6][1] , 
        \i16/rx_fifo/buff[6][2] , \i16/rx_fifo/buff[6][3] , \i16/rx_fifo/buff[6][4] , 
        \i16/rx_fifo/buff[6][5] , \i16/rx_fifo/buff[6][6] , \i16/rx_fifo/buff[6][7] , 
        \i16/rx_fifo/buff[7][0] , \i16/rx_fifo/buff[7][1] , \i16/rx_fifo/buff[7][2] , 
        \i16/rx_fifo/buff[7][3] , \i16/rx_fifo/buff[7][4] , \i16/rx_fifo/buff[7][5] , 
        \i16/rx_fifo/buff[7][6] , \i16/rx_fifo/buff[7][7] , \i16/rx_fifo/buff[8][0] , 
        \i16/rx_fifo/buff[8][1] , \i16/rx_fifo/buff[8][2] , \i16/rx_fifo/buff[8][3] , 
        \i16/rx_fifo/buff[8][4] , \i16/rx_fifo/buff[8][5] , \i16/rx_fifo/buff[8][6] , 
        \i16/rx_fifo/buff[8][7] , \i16/rx_fifo/buff[9][0] , \i16/rx_fifo/buff[9][1] , 
        \i16/rx_fifo/buff[9][2] , \i16/rx_fifo/buff[9][3] , \i16/rx_fifo/buff[9][4] , 
        \i16/rx_fifo/buff[9][5] , \i16/rx_fifo/buff[9][6] , \i16/rx_fifo/buff[9][7] , 
        \i16/rx_fifo/buff[10][0] , \i16/rx_fifo/buff[10][1] , \i16/rx_fifo/buff[10][2] , 
        \i16/rx_fifo/buff[10][3] , \i16/rx_fifo/buff[10][4] , \i16/rx_fifo/buff[10][5] , 
        \i16/rx_fifo/buff[10][6] , \i16/rx_fifo/buff[10][7] , \i16/rx_fifo/buff[11][0] , 
        \i16/rx_fifo/buff[11][1] , \i16/rx_fifo/buff[11][2] , \i16/rx_fifo/buff[11][3] , 
        \i16/rx_fifo/buff[11][4] , \i16/rx_fifo/buff[11][5] , \i16/rx_fifo/buff[11][6] , 
        \i16/rx_fifo/buff[11][7] , \i16/rx_fifo/buff[12][0] , \i16/rx_fifo/buff[12][1] , 
        \i16/rx_fifo/buff[12][2] , \i16/rx_fifo/buff[12][3] , \i16/rx_fifo/buff[12][4] , 
        \i16/rx_fifo/buff[12][5] , \i16/rx_fifo/buff[12][6] , \i16/rx_fifo/buff[12][7] , 
        \i16/rx_fifo/buff[13][0] , \i16/rx_fifo/buff[13][1] , \i16/rx_fifo/buff[13][2] , 
        \i16/rx_fifo/buff[13][3] , \i16/rx_fifo/buff[13][4] , \i16/rx_fifo/buff[13][5] , 
        \i16/rx_fifo/buff[13][6] , \i16/rx_fifo/buff[13][7] , \i16/rx_fifo/buff[14][0] , 
        \i16/rx_fifo/buff[14][1] , \i16/rx_fifo/buff[14][2] , \i16/rx_fifo/buff[14][3] , 
        \i16/rx_fifo/buff[14][4] , \i16/rx_fifo/buff[14][5] , \i16/rx_fifo/buff[14][6] , 
        \i16/rx_fifo/buff[14][7] , \i16/rx_fifo/buff[15][0] , \i16/rx_fifo/buff[15][1] , 
        \i16/rx_fifo/buff[15][2] , \i16/rx_fifo/buff[15][3] , \i16/rx_fifo/buff[15][4] , 
        \i16/rx_fifo/buff[15][5] , \i16/rx_fifo/buff[15][6] , \i16/rx_fifo/buff[15][7] , 
        \i16/rx_fifo/buff[16][0] , \i16/rx_fifo/buff[16][1] , \i16/rx_fifo/buff[16][2] , 
        \i16/rx_fifo/buff[16][3] , \i16/rx_fifo/buff[16][4] , \i16/rx_fifo/buff[16][5] , 
        \i16/rx_fifo/buff[16][6] , \i16/rx_fifo/buff[16][7] , \i16/rx_fifo/buff[17][0] , 
        \i16/rx_fifo/buff[17][1] , \i16/rx_fifo/buff[17][2] , \i16/rx_fifo/buff[17][3] , 
        \i16/rx_fifo/buff[17][4] , \i16/rx_fifo/buff[17][5] , \i16/rx_fifo/buff[17][6] , 
        \i16/rx_fifo/buff[17][7] , \i16/rx_fifo/buff[18][0] , \i16/rx_fifo/buff[18][1] , 
        \i16/rx_fifo/buff[18][2] , \i16/rx_fifo/buff[18][3] , \i16/rx_fifo/buff[18][4] , 
        \i16/rx_fifo/buff[18][5] , \i16/rx_fifo/buff[18][6] , \i16/rx_fifo/buff[18][7] , 
        \i16/rx_fifo/buff[19][0] , \i16/rx_fifo/buff[19][1] , \i16/rx_fifo/buff[19][2] , 
        \i16/rx_fifo/buff[19][3] , \i16/rx_fifo/buff[19][4] , \i16/rx_fifo/buff[19][5] , 
        \i16/rx_fifo/buff[19][6] , \i16/rx_fifo/buff[19][7] , \i16/rx_fifo/buff[20][0] , 
        \i16/rx_fifo/buff[20][1] , \i16/rx_fifo/buff[20][2] , \i16/rx_fifo/buff[20][3] , 
        \i16/rx_fifo/buff[20][4] , \i16/rx_fifo/buff[20][5] , \i16/rx_fifo/buff[20][6] , 
        \i16/rx_fifo/buff[20][7] , \i16/rx_fifo/buff[21][0] , \i16/rx_fifo/buff[21][1] , 
        \i16/rx_fifo/buff[21][2] , \i16/rx_fifo/buff[21][3] , \i16/rx_fifo/buff[21][4] , 
        \i16/rx_fifo/buff[21][5] , \i16/rx_fifo/buff[21][6] , \i16/rx_fifo/buff[21][7] , 
        \i16/rx_fifo/buff[22][0] , \i16/rx_fifo/buff[22][1] , \i16/rx_fifo/buff[22][2] , 
        \i16/rx_fifo/buff[22][3] , \i16/rx_fifo/buff[22][4] , \i16/rx_fifo/buff[22][5] , 
        \i16/rx_fifo/buff[22][6] , \i16/rx_fifo/buff[22][7] , \i16/rx_fifo/buff[23][0] , 
        \i16/rx_fifo/buff[23][1] , \i16/rx_fifo/buff[23][2] , \i16/rx_fifo/buff[23][3] , 
        \i16/rx_fifo/buff[23][4] , \i16/rx_fifo/buff[23][5] , \i16/rx_fifo/buff[23][6] , 
        \i16/rx_fifo/buff[23][7] , \i16/rx_fifo/buff[24][0] , \i16/rx_fifo/buff[24][1] , 
        \i16/rx_fifo/buff[24][2] , \i16/rx_fifo/buff[24][3] , \i16/rx_fifo/buff[24][4] , 
        \i16/rx_fifo/buff[24][5] , \i16/rx_fifo/buff[24][6] , \i16/rx_fifo/buff[24][7] , 
        \i16/rx_fifo/buff[25][0] , \i16/rx_fifo/buff[25][1] , \i16/rx_fifo/buff[25][2] , 
        \i16/rx_fifo/buff[25][3] , \i16/rx_fifo/buff[25][4] , \i16/rx_fifo/buff[25][5] , 
        \i16/rx_fifo/buff[25][6] , \i16/rx_fifo/buff[25][7] , \i16/rx_fifo/buff[26][0] , 
        \i16/rx_fifo/buff[26][1] , \i16/rx_fifo/buff[26][2] , \i16/rx_fifo/buff[26][3] , 
        \i16/rx_fifo/buff[26][4] , \i16/rx_fifo/buff[26][5] , \i16/rx_fifo/buff[26][6] , 
        \i16/rx_fifo/buff[26][7] , \i16/rx_fifo/buff[27][0] , \i16/rx_fifo/buff[27][1] , 
        \i16/rx_fifo/buff[27][2] , \i16/rx_fifo/buff[27][3] , \i16/rx_fifo/buff[27][4] , 
        \i16/rx_fifo/buff[27][5] , \i16/rx_fifo/buff[27][6] , \i16/rx_fifo/buff[27][7] , 
        \i16/rx_fifo/buff[28][0] , \i16/rx_fifo/buff[28][1] , \i16/rx_fifo/buff[28][2] , 
        \i16/rx_fifo/buff[28][3] , \i16/rx_fifo/buff[28][4] , \i16/rx_fifo/buff[28][5] , 
        \i16/rx_fifo/buff[28][6] , \i16/rx_fifo/buff[28][7] , \i16/rx_fifo/buff[29][0] , 
        \i16/rx_fifo/buff[29][1] , \i16/rx_fifo/buff[29][2] , \i16/rx_fifo/buff[29][3] , 
        \i16/rx_fifo/buff[29][4] , \i16/rx_fifo/buff[29][5] , \i16/rx_fifo/buff[29][6] , 
        \i16/rx_fifo/buff[29][7] , \i16/rx_fifo/buff[30][0] , \i16/rx_fifo/buff[30][1] , 
        \i16/rx_fifo/buff[30][2] , \i16/rx_fifo/buff[30][3] , \i16/rx_fifo/buff[30][4] , 
        \i16/rx_fifo/buff[30][5] , \i16/rx_fifo/buff[30][6] , \i16/rx_fifo/buff[30][7] , 
        \i16/rx_fifo/buff[31][0] , \i16/rx_fifo/buff[31][1] , \i16/rx_fifo/buff[31][2] , 
        \i16/rx_fifo/buff[31][3] , \i16/rx_fifo/buff[31][4] , \i16/rx_fifo/buff[31][5] , 
        \i16/rx_fifo/buff[31][6] , \i16/rx_fifo/buff[31][7] , \i16/rx_fifo/buff[32][0] , 
        \i16/rx_fifo/buff[32][1] , \i16/rx_fifo/buff[32][2] , \i16/rx_fifo/buff[32][3] , 
        \i16/rx_fifo/buff[32][4] , \i16/rx_fifo/buff[32][5] , \i16/rx_fifo/buff[32][6] , 
        \i16/rx_fifo/buff[32][7] , \i16/rx_fifo/buff[33][0] , \i16/rx_fifo/buff[33][1] , 
        \i16/rx_fifo/buff[33][2] , \i16/rx_fifo/buff[33][3] , \i16/rx_fifo/buff[33][4] , 
        \i16/rx_fifo/buff[33][5] , \i16/rx_fifo/buff[33][6] , \i16/rx_fifo/buff[33][7] , 
        \i16/rx_fifo/buff[34][0] , \i16/rx_fifo/buff[34][1] , \i16/rx_fifo/buff[34][2] , 
        \i16/rx_fifo/buff[34][3] , \i16/rx_fifo/buff[34][4] , \i16/rx_fifo/buff[34][5] , 
        \i16/rx_fifo/buff[34][6] , \i16/rx_fifo/buff[34][7] , \i16/rx_fifo/buff[35][0] , 
        \i16/rx_fifo/buff[35][1] , \i16/rx_fifo/buff[35][2] , \i16/rx_fifo/buff[35][3] , 
        \i16/rx_fifo/buff[35][4] , \i16/rx_fifo/buff[35][5] , \i16/rx_fifo/buff[35][6] , 
        \i16/rx_fifo/buff[35][7] , \i16/rx_fifo/buff[36][0] , \i16/rx_fifo/buff[36][1] , 
        \i16/rx_fifo/buff[36][2] , \i16/rx_fifo/buff[36][3] , \i16/rx_fifo/buff[36][4] , 
        \i16/rx_fifo/buff[36][5] , \i16/rx_fifo/buff[36][6] , \i16/rx_fifo/buff[36][7] , 
        \i16/rx_fifo/buff[37][0] , \i16/rx_fifo/buff[37][1] , \i16/rx_fifo/buff[37][2] , 
        \i16/rx_fifo/buff[37][3] , \i16/rx_fifo/buff[37][4] , \i16/rx_fifo/buff[37][5] , 
        \i16/rx_fifo/buff[37][6] , \i16/rx_fifo/buff[37][7] , \i16/rx_fifo/buff[38][0] , 
        \i16/rx_fifo/buff[38][1] , \i16/rx_fifo/buff[38][2] , \i16/rx_fifo/buff[38][3] , 
        \i16/rx_fifo/buff[38][4] , \i16/rx_fifo/buff[38][5] , \i16/rx_fifo/buff[38][6] , 
        \i16/rx_fifo/buff[38][7] , \i16/rx_fifo/buff[39][0] , \i16/rx_fifo/buff[39][1] , 
        \i16/rx_fifo/buff[39][2] , \i16/rx_fifo/buff[39][3] , \i16/rx_fifo/buff[39][4] , 
        \i16/rx_fifo/buff[39][5] , \i16/rx_fifo/buff[39][6] , \i16/rx_fifo/buff[39][7] , 
        \i16/rx_fifo/buff[40][0] , \i16/rx_fifo/buff[40][1] , \i16/rx_fifo/buff[40][2] , 
        \i16/rx_fifo/buff[40][3] , \i16/rx_fifo/buff[40][4] , \i16/rx_fifo/buff[40][5] , 
        \i16/rx_fifo/buff[40][6] , \i16/rx_fifo/buff[40][7] , \i16/rx_fifo/buff[41][0] , 
        \i16/rx_fifo/buff[41][1] , \i16/rx_fifo/buff[41][2] , \i16/rx_fifo/buff[41][3] , 
        \i16/rx_fifo/buff[41][4] , \i16/rx_fifo/buff[41][5] , \i16/rx_fifo/buff[41][6] , 
        \i16/rx_fifo/buff[41][7] , \i16/rx_fifo/buff[42][0] , \i16/rx_fifo/buff[42][1] , 
        \i16/rx_fifo/buff[42][2] , \i16/rx_fifo/buff[42][3] , \i16/rx_fifo/buff[42][4] , 
        \i16/rx_fifo/buff[42][5] , \i16/rx_fifo/buff[42][6] , \i16/rx_fifo/buff[42][7] , 
        \i16/rx_fifo/buff[43][0] , \i16/rx_fifo/buff[43][1] , \i16/rx_fifo/buff[43][2] , 
        \i16/rx_fifo/buff[43][3] , \i16/rx_fifo/buff[43][4] , \i16/rx_fifo/buff[43][5] , 
        \i16/rx_fifo/buff[43][6] , \i16/rx_fifo/buff[43][7] , \i16/rx_fifo/buff[44][0] , 
        \i16/rx_fifo/buff[44][1] , \i16/rx_fifo/buff[44][2] , \i16/rx_fifo/buff[44][3] , 
        \i16/rx_fifo/buff[44][4] , \i16/rx_fifo/buff[44][5] , \i16/rx_fifo/buff[44][6] , 
        \i16/rx_fifo/buff[44][7] , \i16/rx_fifo/buff[45][0] , \i16/rx_fifo/buff[45][1] , 
        \i16/rx_fifo/buff[45][2] , \i16/rx_fifo/buff[45][3] , \i16/rx_fifo/buff[45][4] , 
        \i16/rx_fifo/buff[45][5] , \i16/rx_fifo/buff[45][6] , \i16/rx_fifo/buff[45][7] , 
        \i16/rx_fifo/buff[46][0] , \i16/rx_fifo/buff[46][1] , \i16/rx_fifo/buff[46][2] , 
        \i16/rx_fifo/buff[46][3] , \i16/rx_fifo/buff[46][4] , \i16/rx_fifo/buff[46][5] , 
        \i16/rx_fifo/buff[46][6] , \i16/rx_fifo/buff[46][7] , \i16/rx_fifo/buff[47][0] , 
        \i16/rx_fifo/buff[47][1] , \i16/rx_fifo/buff[47][2] , \i16/rx_fifo/buff[47][3] , 
        \i16/rx_fifo/buff[47][4] , \i16/rx_fifo/buff[47][5] , \i16/rx_fifo/buff[47][6] , 
        \i16/rx_fifo/buff[47][7] , \i16/rx_fifo/buff[48][0] , \i16/rx_fifo/buff[48][1] , 
        \i16/rx_fifo/buff[48][2] , \i16/rx_fifo/buff[48][3] , \i16/rx_fifo/buff[48][4] , 
        \i16/rx_fifo/buff[48][5] , \i16/rx_fifo/buff[48][6] , \i16/rx_fifo/buff[48][7] , 
        \i16/rx_fifo/buff[49][0] , \i16/rx_fifo/buff[49][1] , \i16/rx_fifo/buff[49][2] , 
        \i16/rx_fifo/buff[49][3] , \i16/rx_fifo/buff[49][4] , \i16/rx_fifo/buff[49][5] , 
        \i16/rx_fifo/buff[49][6] , \i16/rx_fifo/buff[49][7] , \i16/rx_fifo/buff[50][0] , 
        \i16/rx_fifo/buff[50][1] , \i16/rx_fifo/buff[50][2] , \i16/rx_fifo/buff[50][3] , 
        \i16/rx_fifo/buff[50][4] , \i16/rx_fifo/buff[50][5] , \i16/rx_fifo/buff[50][6] , 
        \i16/rx_fifo/buff[50][7] , \i16/rx_fifo/buff[51][0] , \i16/rx_fifo/buff[51][1] , 
        \i16/rx_fifo/buff[51][2] , \i16/rx_fifo/buff[51][3] , \i16/rx_fifo/buff[51][4] , 
        \i16/rx_fifo/buff[51][5] , \i16/rx_fifo/buff[51][6] , \i16/rx_fifo/buff[51][7] , 
        \i16/rx_fifo/buff[52][0] , \i16/rx_fifo/buff[52][1] , \i16/rx_fifo/buff[52][2] , 
        \i16/rx_fifo/buff[52][3] , \i16/rx_fifo/buff[52][4] , \i16/rx_fifo/buff[52][5] , 
        \i16/rx_fifo/buff[52][6] , \i16/rx_fifo/buff[52][7] , \i16/rx_fifo/buff[53][0] , 
        \i16/rx_fifo/buff[53][1] , \i16/rx_fifo/buff[53][2] , \i16/rx_fifo/buff[53][3] , 
        \i16/rx_fifo/buff[53][4] , \i16/rx_fifo/buff[53][5] , \i16/rx_fifo/buff[53][6] , 
        \i16/rx_fifo/buff[53][7] , \i16/rx_fifo/buff[54][0] , \i16/rx_fifo/buff[54][1] , 
        \i16/rx_fifo/buff[54][2] , \i16/rx_fifo/buff[54][3] , \i16/rx_fifo/buff[54][4] , 
        \i16/rx_fifo/buff[54][5] , \i16/rx_fifo/buff[54][6] , \i16/rx_fifo/buff[54][7] , 
        \i16/rx_fifo/buff[55][0] , \i16/rx_fifo/buff[55][1] , \i16/rx_fifo/buff[55][2] , 
        \i16/rx_fifo/buff[55][3] , \i16/rx_fifo/buff[55][4] , \i16/rx_fifo/buff[55][5] , 
        \i16/rx_fifo/buff[55][6] , \i16/rx_fifo/buff[55][7] , \i16/rx_fifo/buff[56][0] , 
        \i16/rx_fifo/buff[56][1] , \i16/rx_fifo/buff[56][2] , \i16/rx_fifo/buff[56][3] , 
        \i16/rx_fifo/buff[56][4] , \i16/rx_fifo/buff[56][5] , \i16/rx_fifo/buff[56][6] , 
        \i16/rx_fifo/buff[56][7] , \i16/rx_fifo/buff[57][0] , \i16/rx_fifo/buff[57][1] , 
        \i16/rx_fifo/buff[57][2] , \i16/rx_fifo/buff[57][3] , \i16/rx_fifo/buff[57][4] , 
        \i16/rx_fifo/buff[57][5] , \i16/rx_fifo/buff[57][6] , \i16/rx_fifo/buff[57][7] , 
        \i16/rx_fifo/buff[58][0] , \i16/rx_fifo/buff[58][1] , \i16/rx_fifo/buff[58][2] , 
        \i16/rx_fifo/buff[58][3] , \i16/rx_fifo/buff[58][4] , \i16/rx_fifo/buff[58][5] , 
        \i16/rx_fifo/buff[58][6] , \i16/rx_fifo/buff[58][7] , \i16/rx_fifo/buff[59][0] , 
        \i16/rx_fifo/buff[59][1] , \i16/rx_fifo/buff[59][2] , \i16/rx_fifo/buff[59][3] , 
        \i16/rx_fifo/buff[59][4] , \i16/rx_fifo/buff[59][5] , \i16/rx_fifo/buff[59][6] , 
        \i16/rx_fifo/buff[59][7] , \i16/rx_fifo/buff[60][0] , \i16/rx_fifo/buff[60][1] , 
        \i16/rx_fifo/buff[60][2] , \i16/rx_fifo/buff[60][3] , \i16/rx_fifo/buff[60][4] , 
        \i16/rx_fifo/buff[60][5] , \i16/rx_fifo/buff[60][6] , \i16/rx_fifo/buff[60][7] , 
        \i16/rx_fifo/buff[61][0] , \i16/rx_fifo/buff[61][1] , \i16/rx_fifo/buff[61][2] , 
        \i16/rx_fifo/buff[61][3] , \i16/rx_fifo/buff[61][4] , \i16/rx_fifo/buff[61][5] , 
        \i16/rx_fifo/buff[61][6] , \i16/rx_fifo/buff[61][7] , \i16/rx_fifo/buff[62][0] , 
        \i16/rx_fifo/buff[62][1] , \i16/rx_fifo/buff[62][2] , \i16/rx_fifo/buff[62][3] , 
        \i16/rx_fifo/buff[62][4] , \i16/rx_fifo/buff[62][5] , \i16/rx_fifo/buff[62][6] , 
        \i16/rx_fifo/buff[62][7] , \i16/rx_fifo/buff[63][0] , \i16/rx_fifo/buff[63][1] , 
        \i16/rx_fifo/buff[63][2] , \i16/rx_fifo/buff[63][3] , \i16/rx_fifo/buff[63][4] , 
        \i16/rx_fifo/buff[63][5] , \i16/rx_fifo/buff[63][6] , \i16/rx_fifo/buff[63][7] , 
        \i16/rx_fifo/buff[64][0] , \i16/rx_fifo/buff[64][1] , \i16/rx_fifo/buff[64][2] , 
        \i16/rx_fifo/buff[64][3] , \i16/rx_fifo/buff[64][4] , \i16/rx_fifo/buff[64][5] , 
        \i16/rx_fifo/buff[64][6] , \i16/rx_fifo/buff[64][7] , \i16/rx_fifo/buff[65][0] , 
        \i16/rx_fifo/buff[65][1] , \i16/rx_fifo/buff[65][2] , \i16/rx_fifo/buff[65][3] , 
        \i16/rx_fifo/buff[65][4] , \i16/rx_fifo/buff[65][5] , \i16/rx_fifo/buff[65][6] , 
        \i16/rx_fifo/buff[65][7] , \i16/rx_fifo/buff[66][0] , \i16/rx_fifo/buff[66][1] , 
        \i16/rx_fifo/buff[66][2] , \i16/rx_fifo/buff[66][3] , \i16/rx_fifo/buff[66][4] , 
        \i16/rx_fifo/buff[66][5] , \i16/rx_fifo/buff[66][6] , \i16/rx_fifo/buff[66][7] , 
        \i16/rx_fifo/buff[67][0] , \i16/rx_fifo/buff[67][1] , \i16/rx_fifo/buff[67][2] , 
        \i16/rx_fifo/buff[67][3] , \i16/rx_fifo/buff[67][4] , \i16/rx_fifo/buff[67][5] , 
        \i16/rx_fifo/buff[67][6] , \i16/rx_fifo/buff[67][7] , \i16/rx_fifo/buff[68][0] , 
        \i16/rx_fifo/buff[68][1] , \i16/rx_fifo/buff[68][2] , \i16/rx_fifo/buff[68][3] , 
        \i16/rx_fifo/buff[68][4] , \i16/rx_fifo/buff[68][5] , \i16/rx_fifo/buff[68][6] , 
        \i16/rx_fifo/buff[68][7] , \i16/rx_fifo/buff[69][0] , \i16/rx_fifo/buff[69][1] , 
        \i16/rx_fifo/buff[69][2] , \i16/rx_fifo/buff[69][3] , \i16/rx_fifo/buff[69][4] , 
        \i16/rx_fifo/buff[69][5] , \i16/rx_fifo/buff[69][6] , \i16/rx_fifo/buff[69][7] , 
        \i16/rx_fifo/buff[70][0] , \i16/rx_fifo/buff[70][1] , \i16/rx_fifo/buff[70][2] , 
        \i16/rx_fifo/buff[70][3] , \i16/rx_fifo/buff[70][4] , \i16/rx_fifo/buff[70][5] , 
        \i16/rx_fifo/buff[70][6] , \i16/rx_fifo/buff[70][7] , \i16/rx_fifo/buff[71][0] , 
        \i16/rx_fifo/buff[71][1] , \i16/rx_fifo/buff[71][2] , \i16/rx_fifo/buff[71][3] , 
        \i16/rx_fifo/buff[71][4] , \i16/rx_fifo/buff[71][5] , \i16/rx_fifo/buff[71][6] , 
        \i16/rx_fifo/buff[71][7] , \i16/rx_fifo/buff[72][0] , \i16/rx_fifo/buff[72][1] , 
        \i16/rx_fifo/buff[72][2] , \i16/rx_fifo/buff[72][3] , \i16/rx_fifo/buff[72][4] , 
        \i16/rx_fifo/buff[72][5] , \i16/rx_fifo/buff[72][6] , \i16/rx_fifo/buff[72][7] , 
        \i16/rx_fifo/buff[73][0] , \i16/rx_fifo/buff[73][1] , \i16/rx_fifo/buff[73][2] , 
        \i16/rx_fifo/buff[73][3] , \i16/rx_fifo/buff[73][4] , \i16/rx_fifo/buff[73][5] , 
        \i16/rx_fifo/buff[73][6] , \i16/rx_fifo/buff[73][7] , \i16/rx_fifo/buff[74][0] , 
        \i16/rx_fifo/buff[74][1] , \i16/rx_fifo/buff[74][2] , \i16/rx_fifo/buff[74][3] , 
        \i16/rx_fifo/buff[74][4] , \i16/rx_fifo/buff[74][5] , \i16/rx_fifo/buff[74][6] , 
        \i16/rx_fifo/buff[74][7] , \i16/rx_fifo/buff[75][0] , \i16/rx_fifo/buff[75][1] , 
        \i16/rx_fifo/buff[75][2] , \i16/rx_fifo/buff[75][3] , \i16/rx_fifo/buff[75][4] , 
        \i16/rx_fifo/buff[75][5] , \i16/rx_fifo/buff[75][6] , \i16/rx_fifo/buff[75][7] , 
        \i16/rx_fifo/buff[76][0] , \i16/rx_fifo/buff[76][1] , \i16/rx_fifo/buff[76][2] , 
        \i16/rx_fifo/buff[76][3] , \i16/rx_fifo/buff[76][4] , \i16/rx_fifo/buff[76][5] , 
        \i16/rx_fifo/buff[76][6] , \i16/rx_fifo/buff[76][7] , \i16/rx_fifo/buff[77][0] , 
        \i16/rx_fifo/buff[77][1] , \i16/rx_fifo/buff[77][2] , \i16/rx_fifo/buff[77][3] , 
        \i16/rx_fifo/buff[77][4] , \i16/rx_fifo/buff[77][5] , \i16/rx_fifo/buff[77][6] , 
        \i16/rx_fifo/buff[77][7] , \i16/rx_fifo/buff[78][0] , \i16/rx_fifo/buff[78][1] , 
        \i16/rx_fifo/buff[78][2] , \i16/rx_fifo/buff[78][3] , \i16/rx_fifo/buff[78][4] , 
        \i16/rx_fifo/buff[78][5] , \i16/rx_fifo/buff[78][6] , \i16/rx_fifo/buff[78][7] , 
        \i16/rx_fifo/buff[79][0] , \i16/rx_fifo/buff[79][1] , \i16/rx_fifo/buff[79][2] , 
        \i16/rx_fifo/buff[79][3] , \i16/rx_fifo/buff[79][4] , \i16/rx_fifo/buff[79][5] , 
        \i16/rx_fifo/buff[79][6] , \i16/rx_fifo/buff[79][7] , \i16/rx_fifo/buff[80][0] , 
        \i16/rx_fifo/buff[80][1] , \i16/rx_fifo/buff[80][2] , \i16/rx_fifo/buff[80][3] , 
        \i16/rx_fifo/buff[80][4] , \i16/rx_fifo/buff[80][5] , \i16/rx_fifo/buff[80][6] , 
        \i16/rx_fifo/buff[80][7] , \i16/rx_fifo/buff[81][0] , \i16/rx_fifo/buff[81][1] , 
        \i16/rx_fifo/buff[81][2] , \i16/rx_fifo/buff[81][3] , \i16/rx_fifo/buff[81][4] , 
        \i16/rx_fifo/buff[81][5] , \i16/rx_fifo/buff[81][6] , \i16/rx_fifo/buff[81][7] , 
        \i16/rx_fifo/buff[82][0] , \i16/rx_fifo/buff[82][1] , \i16/rx_fifo/buff[82][2] , 
        \i16/rx_fifo/buff[82][3] , \i16/rx_fifo/buff[82][4] , \i16/rx_fifo/buff[82][5] , 
        \i16/rx_fifo/buff[82][6] , \i16/rx_fifo/buff[82][7] , \i16/rx_fifo/buff[83][0] , 
        \i16/rx_fifo/buff[83][1] , \i16/rx_fifo/buff[83][2] , \i16/rx_fifo/buff[83][3] , 
        \i16/rx_fifo/buff[83][4] , \i16/rx_fifo/buff[83][5] , \i16/rx_fifo/buff[83][6] , 
        \i16/rx_fifo/buff[83][7] , \i16/rx_fifo/buff[84][0] , \i16/rx_fifo/buff[84][1] , 
        \i16/rx_fifo/buff[84][2] , \i16/rx_fifo/buff[84][3] , \i16/rx_fifo/buff[84][4] , 
        \i16/rx_fifo/buff[84][5] , \i16/rx_fifo/buff[84][6] , \i16/rx_fifo/buff[84][7] , 
        \i16/rx_fifo/buff[85][0] , \i16/rx_fifo/buff[85][1] , \i16/rx_fifo/buff[85][2] , 
        \i16/rx_fifo/buff[85][3] , \i16/rx_fifo/buff[85][4] , \i16/rx_fifo/buff[85][5] , 
        \i16/rx_fifo/buff[85][6] , \i16/rx_fifo/buff[85][7] , \i16/rx_fifo/buff[86][0] , 
        \i16/rx_fifo/buff[86][1] , \i16/rx_fifo/buff[86][2] , \i16/rx_fifo/buff[86][3] , 
        \i16/rx_fifo/buff[86][4] , \i16/rx_fifo/buff[86][5] , \i16/rx_fifo/buff[86][6] , 
        \i16/rx_fifo/buff[86][7] , \i16/rx_fifo/buff[87][0] , \i16/rx_fifo/buff[87][1] , 
        \i16/rx_fifo/buff[87][2] , \i16/rx_fifo/buff[87][3] , \i16/rx_fifo/buff[87][4] , 
        \i16/rx_fifo/buff[87][5] , \i16/rx_fifo/buff[87][6] , \i16/rx_fifo/buff[87][7] , 
        \i16/rx_fifo/buff[88][0] , \i16/rx_fifo/buff[88][1] , \i16/rx_fifo/buff[88][2] , 
        \i16/rx_fifo/buff[88][3] , \i16/rx_fifo/buff[88][4] , \i16/rx_fifo/buff[88][5] , 
        \i16/rx_fifo/buff[88][6] , \i16/rx_fifo/buff[88][7] , \i16/rx_fifo/buff[89][0] , 
        \i16/rx_fifo/buff[89][1] , \i16/rx_fifo/buff[89][2] , \i16/rx_fifo/buff[89][3] , 
        \i16/rx_fifo/buff[89][4] , \i16/rx_fifo/buff[89][5] , \i16/rx_fifo/buff[89][6] , 
        \i16/rx_fifo/buff[89][7] , \i16/rx_fifo/buff[90][0] , \i16/rx_fifo/buff[90][1] , 
        \i16/rx_fifo/buff[90][2] , \i16/rx_fifo/buff[90][3] , \i16/rx_fifo/buff[90][4] , 
        \i16/rx_fifo/buff[90][5] , \i16/rx_fifo/buff[90][6] , \i16/rx_fifo/buff[90][7] , 
        \i16/rx_fifo/buff[91][0] , \i16/rx_fifo/buff[91][1] , \i16/rx_fifo/buff[91][2] , 
        \i16/rx_fifo/buff[91][3] , \i16/rx_fifo/buff[91][4] , \i16/rx_fifo/buff[91][5] , 
        \i16/rx_fifo/buff[91][6] , \i16/rx_fifo/buff[91][7] , \i16/rx_fifo/buff[92][0] , 
        \i16/rx_fifo/buff[92][1] , \i16/rx_fifo/buff[92][2] , \i16/rx_fifo/buff[92][3] , 
        \i16/rx_fifo/buff[92][4] , \i16/rx_fifo/buff[92][5] , \i16/rx_fifo/buff[92][6] , 
        \i16/rx_fifo/buff[92][7] , \i16/rx_fifo/buff[93][0] , \i16/rx_fifo/buff[93][1] , 
        \i16/rx_fifo/buff[93][2] , \i16/rx_fifo/buff[93][3] , \i16/rx_fifo/buff[93][4] , 
        \i16/rx_fifo/buff[93][5] , \i16/rx_fifo/buff[93][6] , \i16/rx_fifo/buff[93][7] , 
        \i16/rx_fifo/buff[94][0] , \i16/rx_fifo/buff[94][1] , \i16/rx_fifo/buff[94][2] , 
        \i16/rx_fifo/buff[94][3] , \i16/rx_fifo/buff[94][4] , \i16/rx_fifo/buff[94][5] , 
        \i16/rx_fifo/buff[94][6] , \i16/rx_fifo/buff[94][7] , \i16/rx_fifo/buff[95][0] , 
        \i16/rx_fifo/buff[95][1] , \i16/rx_fifo/buff[95][2] , \i16/rx_fifo/buff[95][3] , 
        \i16/rx_fifo/buff[95][4] , \i16/rx_fifo/buff[95][5] , \i16/rx_fifo/buff[95][6] , 
        \i16/rx_fifo/buff[95][7] , \i16/rx_fifo/buff[96][0] , \i16/rx_fifo/buff[96][1] , 
        \i16/rx_fifo/buff[96][2] , \i16/rx_fifo/buff[96][3] , \i16/rx_fifo/buff[96][4] , 
        \i16/rx_fifo/buff[96][5] , \i16/rx_fifo/buff[96][6] , \i16/rx_fifo/buff[96][7] , 
        \i16/rx_fifo/buff[97][0] , \i16/rx_fifo/buff[97][1] , \i16/rx_fifo/buff[97][2] , 
        \i16/rx_fifo/buff[97][3] , \i16/rx_fifo/buff[97][4] , \i16/rx_fifo/buff[97][5] , 
        \i16/rx_fifo/buff[97][6] , \i16/rx_fifo/buff[97][7] , \i16/rx_fifo/buff[98][0] , 
        \i16/rx_fifo/buff[98][1] , \i16/rx_fifo/buff[98][2] , \i16/rx_fifo/buff[98][3] , 
        \i16/rx_fifo/buff[98][4] , \i16/rx_fifo/buff[98][5] , \i16/rx_fifo/buff[98][6] , 
        \i16/rx_fifo/buff[98][7] , \i16/rx_fifo/buff[99][0] , \i16/rx_fifo/buff[99][1] , 
        \i16/rx_fifo/buff[99][2] , \i16/rx_fifo/buff[99][3] , \i16/rx_fifo/buff[99][4] , 
        \i16/rx_fifo/buff[99][5] , \i16/rx_fifo/buff[99][6] , \i16/rx_fifo/buff[99][7] , 
        \i16/rx_fifo/buff[100][0] , \i16/rx_fifo/buff[100][1] , \i16/rx_fifo/buff[100][2] , 
        \i16/rx_fifo/buff[100][3] , \i16/rx_fifo/buff[100][4] , \i16/rx_fifo/buff[100][5] , 
        \i16/rx_fifo/buff[100][6] , \i16/rx_fifo/buff[100][7] , \i16/rx_fifo/buff[101][0] , 
        \i16/rx_fifo/buff[101][1] , \i16/rx_fifo/buff[101][2] , \i16/rx_fifo/buff[101][3] , 
        \i16/rx_fifo/buff[101][4] , \i16/rx_fifo/buff[101][5] , \i16/rx_fifo/buff[101][6] , 
        \i16/rx_fifo/buff[101][7] , \i16/rx_fifo/buff[102][0] , \i16/rx_fifo/buff[102][1] , 
        \i16/rx_fifo/buff[102][2] , \i16/rx_fifo/buff[102][3] , \i16/rx_fifo/buff[102][4] , 
        \i16/rx_fifo/buff[102][5] , \i16/rx_fifo/buff[102][6] , \i16/rx_fifo/buff[102][7] , 
        \i16/rx_fifo/buff[103][0] , \i16/rx_fifo/buff[103][1] , \i16/rx_fifo/buff[103][2] , 
        \i16/rx_fifo/buff[103][3] , \i16/rx_fifo/buff[103][4] , \i16/rx_fifo/buff[103][5] , 
        \i16/rx_fifo/buff[103][6] , \i16/rx_fifo/buff[103][7] , \i16/rx_fifo/buff[104][0] , 
        \i16/rx_fifo/buff[104][1] , \i16/rx_fifo/buff[104][2] , \i16/rx_fifo/buff[104][3] , 
        \i16/rx_fifo/buff[104][4] , \i16/rx_fifo/buff[104][5] , \i16/rx_fifo/buff[104][6] , 
        \i16/rx_fifo/buff[104][7] , \i16/rx_fifo/buff[105][0] , \i16/rx_fifo/buff[105][1] , 
        \i16/rx_fifo/buff[105][2] , \i16/rx_fifo/buff[105][3] , \i16/rx_fifo/buff[105][4] , 
        \i16/rx_fifo/buff[105][5] , \i16/rx_fifo/buff[105][6] , \i16/rx_fifo/buff[105][7] , 
        \i16/rx_fifo/buff[106][0] , \i16/rx_fifo/buff[106][1] , \i16/rx_fifo/buff[106][2] , 
        \i16/rx_fifo/buff[106][3] , \i16/rx_fifo/buff[106][4] , \i16/rx_fifo/buff[106][5] , 
        \i16/rx_fifo/buff[106][6] , \i16/rx_fifo/buff[106][7] , \i16/rx_fifo/buff[107][0] , 
        \i16/rx_fifo/buff[107][1] , \i16/rx_fifo/buff[107][2] , \i16/rx_fifo/buff[107][3] , 
        \i16/rx_fifo/buff[107][4] , \i16/rx_fifo/buff[107][5] , \i16/rx_fifo/buff[107][6] , 
        \i16/rx_fifo/buff[107][7] , \i16/rx_fifo/buff[108][0] , \i16/rx_fifo/buff[108][1] , 
        \i16/rx_fifo/buff[108][2] , \i16/rx_fifo/buff[108][3] , \i16/rx_fifo/buff[108][4] , 
        \i16/rx_fifo/buff[108][5] , \i16/rx_fifo/buff[108][6] , \i16/rx_fifo/buff[108][7] , 
        \i16/rx_fifo/buff[109][0] , \i16/rx_fifo/buff[109][1] , \i16/rx_fifo/buff[109][2] , 
        \i16/rx_fifo/buff[109][3] , \i16/rx_fifo/buff[109][4] , n3179, 
        \i16/rx_fifo/buff[109][5] , \i16/rx_fifo/buff[109][6] , n3182, 
        n3183, \i16/rx_fifo/buff[109][7] , n3185, n3186, \i16/rx_fifo/buff[110][0] , 
        \i16/rx_fifo/buff[110][1] , n3189, n3190, \i16/rx_fifo/buff[110][2] , 
        n3192, n3193, \i16/rx_fifo/buff[110][3] , \i16/rx_fifo/buff[110][4] , 
        n3196, n3197, \i16/rx_fifo/buff[110][5] , \i16/rx_fifo/buff[110][6] , 
        \i16/rx_fifo/buff[110][7] , \i16/rx_fifo/buff[111][0] , n3202, 
        \i16/rx_fifo/buff[111][1] , \i16/rx_fifo/buff[111][2] , n3205, 
        n3206, \i16/rx_fifo/buff[111][3] , n3208, n3209, \i16/rx_fifo/buff[111][4] , 
        \i16/rx_fifo/buff[111][5] , n3212, n3213, \i16/rx_fifo/buff[111][6] , 
        n3215, n3216, \i16/rx_fifo/buff[111][7] , \i16/rx_fifo/buff[112][0] , 
        n3219, n3220, \i16/rx_fifo/buff[112][1] , \i16/rx_fifo/buff[112][2] , 
        \i16/rx_fifo/buff[112][3] , \i16/rx_fifo/buff[112][4] , \i16/rx_fifo/buff[112][5] , 
        n3226, \i16/rx_fifo/buff[112][6] , n3228, n3229, \i16/rx_fifo/buff[112][7] , 
        n3231, n3232, \i16/rx_fifo/buff[113][0] , n3234, n3235, \i16/rx_fifo/buff[113][1] , 
        n3237, n3238, \i16/rx_fifo/buff[113][2] , \i16/rx_fifo/buff[113][3] , 
        \i16/rx_fifo/buff[113][4] , \i16/rx_fifo/buff[113][5] , \i16/rx_fifo/buff[113][6] , 
        \i16/rx_fifo/buff[113][7] , \i16/rx_fifo/buff[114][0] , \i16/rx_fifo/buff[114][1] , 
        \i16/rx_fifo/buff[114][2] , \i16/rx_fifo/buff[114][3] , \i16/rx_fifo/buff[114][4] , 
        \i16/rx_fifo/buff[114][5] , \i16/rx_fifo/buff[114][6] , \i16/rx_fifo/buff[114][7] , 
        \i16/rx_fifo/buff[115][0] , \i16/rx_fifo/buff[115][1] , \i16/rx_fifo/buff[115][2] , 
        \i16/rx_fifo/buff[115][3] , \i16/rx_fifo/buff[115][4] , \i16/rx_fifo/buff[115][5] , 
        \i16/rx_fifo/buff[115][6] , n3260, n3261, \i16/rx_fifo/buff[115][7] , 
        \i16/rx_fifo/buff[116][0] , \i16/rx_fifo/buff[116][1] , \i16/rx_fifo/buff[116][2] , 
        \i16/rx_fifo/buff[116][3] , n3267, \i16/rx_fifo/buff[116][4] , 
        n3269, n3270, \i16/rx_fifo/buff[116][5] , \i16/rx_fifo/buff[116][6] , 
        n3273, n3274, \i16/rx_fifo/buff[116][7] , n3276, \i16/rx_fifo/buff[117][0] , 
        \i16/rx_fifo/buff[117][1] , \i16/rx_fifo/buff[117][2] , \i16/rx_fifo/buff[117][3] , 
        \i16/rx_fifo/buff[117][4] , n3282, \i16/rx_fifo/buff[117][5] , 
        n3284, n3285, \i16/rx_fifo/buff[117][6] , \i16/rx_fifo/buff[117][7] , 
        n3288, n3289, \i16/rx_fifo/buff[118][0] , \i16/rx_fifo/buff[118][1] , 
        \i16/rx_fifo/buff[118][2] , \i16/rx_fifo/buff[118][3] , \i16/rx_fifo/buff[118][4] , 
        n3295, \i16/rx_fifo/buff[118][5] , \i16/rx_fifo/buff[118][6] , 
        \i16/rx_fifo/buff[118][7] , \i16/rx_fifo/buff[119][0] , n3300, 
        \i16/rx_fifo/buff[119][1] , n3302, \i16/rx_fifo/buff[119][2] , 
        \i16/rx_fifo/buff[119][3] , \i16/rx_fifo/buff[119][4] , \i16/rx_fifo/buff[119][5] , 
        n3307, \i16/rx_fifo/buff[119][6] , \i16/rx_fifo/buff[119][7] , 
        n3310, n3311, \i16/rx_fifo/buff[120][0] , n3313, n3314, \i16/rx_fifo/buff[120][1] , 
        n3316, n3317, \i16/rx_fifo/buff[120][2] , \i16/rx_fifo/buff[120][3] , 
        \i16/rx_fifo/buff[120][4] , \i16/rx_fifo/buff[120][5] , \i16/rx_fifo/buff[120][6] , 
        \i16/rx_fifo/buff[120][7] , n3324, \i16/rx_fifo/buff[121][0] , 
        n3326, n3327, \i16/rx_fifo/buff[121][1] , n3329, n3330, \i16/rx_fifo/buff[121][2] , 
        \i16/rx_fifo/buff[121][3] , n3333, n3334, \i16/rx_fifo/buff[121][4] , 
        \i16/rx_fifo/buff[121][5] , \i16/rx_fifo/buff[121][6] , \i16/rx_fifo/buff[121][7] , 
        n3339, n3340, \i16/rx_fifo/buff[122][0] , \i16/rx_fifo/buff[122][1] , 
        n3343, n3344, \i16/rx_fifo/buff[122][2] , n3346, n3347, \i16/rx_fifo/buff[122][3] , 
        \i16/rx_fifo/buff[122][4] , n3350, n3351, \i16/rx_fifo/buff[122][5] , 
        \i16/rx_fifo/buff[122][6] , \i16/rx_fifo/buff[122][7] , \i16/rx_fifo/buff[123][0] , 
        \i16/rx_fifo/buff[123][1] , n3357, n3358, \i16/rx_fifo/buff[123][2] , 
        \i16/rx_fifo/buff[123][3] , \i16/rx_fifo/buff[123][4] , n3362, 
        n3363, \i16/rx_fifo/buff[123][5] , \i16/rx_fifo/buff[123][6] , 
        n3366, n3367, \i16/rx_fifo/buff[123][7] , \i16/rx_fifo/buff[124][0] , 
        n3370, n3371, \i16/rx_fifo/buff[124][1] , \i16/rx_fifo/buff[124][2] , 
        \i16/rx_fifo/buff[124][3] , n3375, n3376, \i16/rx_fifo/buff[124][4] , 
        \i16/rx_fifo/buff[124][5] , n3379, n3380, \i16/rx_fifo/buff[124][6] , 
        \i16/rx_fifo/buff[124][7] , \i16/rx_fifo/buff[125][0] , \i16/rx_fifo/buff[125][1] , 
        n3385, n3386, \i16/rx_fifo/buff[125][2] , \i16/rx_fifo/buff[125][3] , 
        n3389, n3390, \i16/rx_fifo/buff[125][4] , n3392, n3393, \i16/rx_fifo/buff[125][5] , 
        \i16/rx_fifo/buff[125][6] , n3396, n3397, \i16/rx_fifo/buff[125][7] , 
        n3399, n3400, \i16/rx_fifo/buff[126][0] , \i16/rx_fifo/buff[126][1] , 
        n3403, n3404, \i16/rx_fifo/buff[126][2] , n3406, n3407, \i16/rx_fifo/buff[126][3] , 
        \i16/rx_fifo/buff[126][4] , n3410, n3411, \i16/rx_fifo/buff[126][5] , 
        \i16/rx_fifo/buff[126][6] , \i16/rx_fifo/buff[126][7] , \i16/rx_fifo/buff[127][0] , 
        n3416, \i16/rx_fifo/buff[127][1] , \i16/rx_fifo/buff[127][2] , 
        n3419, n3420, \i16/rx_fifo/buff[127][3] , n3422, n3423, \i16/rx_fifo/buff[127][4] , 
        \i16/rx_fifo/buff[127][5] , n3426, n3427, \i16/rx_fifo/buff[127][6] , 
        \i16/rx_fifo/buff[127][7] , \spi_slave_inst/n94 , ceg_net49, \spi_slave_inst/n95 , 
        \spi_slave_inst/n56 , ceg_net40, \spi_slave_inst/n57 , \spi_slave_inst/sync_tx_en[0] , 
        \spi_slave_inst/n96 , \spi_slave_inst/n97 , tx_en, \spi_slave_inst/n58 , 
        \spi_slave_inst/sync_mosi[0] , \spi_slave_inst/n73 , ceg_net23, 
        \spi_slave_inst/n98 , \spi_slave_inst/n139 , ceg_net77, ceg_net98, 
        \spi_slave_inst/n68 , ceg_net34, ceg_net37, \spi_slave_inst/n54 , 
        \spi_slave_inst/n93 , \spi_slave_inst/n55 , \spi_slave_inst/n92 , 
        \spi_slave_inst/n138 , \spi_slave_inst/n137 , \spi_slave_inst/n136 , 
        \spi_slave_inst/n135 , \spi_slave_inst/n134 , \spi_slave_inst/n133 , 
        \spi_slave_inst/n132 , \spi_slave_inst/n173 , \spi_slave_inst/n172 , 
        \spi_slave_inst/n171 , \spi_slave_inst/n170 , \spi_slave_inst/n169 , 
        \spi_slave_inst/n168 , \spi_slave_inst/n167 , \led_inst/n41 , 
        \led_inst/n42 , \led_inst/n43 , \led_inst/n44 , \led_inst/n45 , 
        \led_inst/n48 , \led_inst/n46 , \led_inst/n47 , \led_inst/n142 , 
        \data_to_led[0] , rx_en_led, \led_inst/LessThan_21/n48 , \led_inst/n141 , 
        \led_inst/n140 , \led_inst/n139 , \led_inst/n138 , \led_inst/n137 , 
        \led_inst/n136 , \led_inst/n135 , \led_inst/n134 , \led_inst/n133 , 
        \led_inst/n132 , \led_inst/n131 , \led_inst/n130 , \led_inst/n129 , 
        \led_inst/n128 , \led_inst/n127 , \led_inst/n126 , \led_inst/n125 , 
        \led_inst/n124 , \led_inst/n123 , \led_inst/n122 , \led_inst/n121 , 
        \led_inst/n120 , \led_inst/n119 , \data_to_led[1] , \data_to_led[2] , 
        \data_to_led[3] , \data_to_led[4] , \data_to_led[5] , \data_to_led[6] , 
        \data_to_led[7] , \data_to_gpo[0] , rx_en_gpo, \data_to_gpo[1] , 
        \data_to_gpo[2] , \data_to_gpo[3] , \data_to_gpo[4] , \data_to_gpo[5] , 
        \data_to_gpo[6] , \data_to_gpo[7] , \data_to_fifo[2] , \i14/n129 , 
        \data_to_fifo[1] , \data_to_fifo[0] , \data_to_fifo[7] , \i14/n130 , 
        \tx_dac_fsm_inst/n68 , \tx_dac_fsm_inst/n42 , \tx_dac_fsm_inst/n344 , 
        n3556, n3557, \tx_dac_fsm_inst/n67 , \tx_dac_fsm_inst/n66 , 
        \tx_dac_fsm_inst/n65 , n3561, n3562, \data_to_fifo[6] , n3564, 
        n3565, \tx_dac_fsm_inst/n258 , \tx_dac_fsm_inst/n64 , \tx_dac_fsm_inst/n284 , 
        data_to_dac, rx_en_dac, \~tx_dac_fsm_inst/n431 , \~tx_dac_fsm_inst/n436 , 
        \~tx_dac_fsm_inst/n441 , n3583, n3584, n3585, n3586, \tx_dac_fsm_inst/n257 , 
        \tx_dac_fsm_inst/n256 , \tx_dac_fsm_inst/n255 , \tx_dac_fsm_inst/n254 , 
        \tx_dac_fsm_inst/n253 , \tx_dac_fsm_inst/n283 , \tx_dac_fsm_inst/n282 , 
        \tx_dac_fsm_inst/n281 , \tx_dac_fsm_inst/n280 , \tx_dac_fsm_inst/n279 , 
        \fifo_inst/n153 , ceg_net146, \fifo_inst/n162 , ceg_net164, 
        \data_to_fifo_length[0] , rx_en_fifo_length, rx_en_fifo, tx_en_fifo, 
        \fifo_inst/n144 , ceg_net418, \fifo_inst/n152 , \fifo_inst/n151 , 
        \fifo_inst/n150 , \fifo_inst/n149 , \fifo_inst/n148 , \fifo_inst/n147 , 
        \fifo_inst/n146 , \fifo_inst/n161 , \fifo_inst/n160 , \fifo_inst/n159 , 
        \fifo_inst/n158 , \fifo_inst/n157 , \fifo_inst/n156 , \fifo_inst/n155 , 
        \data_to_fifo_length[1] , \data_to_fifo_length[2] , \data_to_fifo_length[3] , 
        \data_to_fifo_length[4] , \data_to_fifo_length[5] , \data_to_fifo_length[6] , 
        \data_to_fifo_length[7] , \i14/n132 , \data_to_fifo[4] , \i14/n131 , 
        \data_to_fifo[5] , \data_to_fifo[3] , \fifo_inst/n143 , \fifo_inst/n142 , 
        \fifo_inst/n141 , \fifo_inst/n140 , \fifo_inst/n139 , \fifo_inst/n138 , 
        \fifo_inst/n137 , \tx_fifo/n153 , ceg_net234, \tx_fifo/n162 , 
        ceg_net252, \data_to_tx_packet_len_reg[0] , rx_en_tx_packet_len, 
        rx_en_tx_packet, tx_en_tx_packet, \tx_fifo/n144 , ceg_net458, 
        \tx_fifo/n152 , \tx_fifo/n151 , \tx_fifo/n150 , \tx_fifo/n149 , 
        \tx_fifo/n148 , \tx_fifo/n147 , \tx_fifo/n146 , \tx_fifo/n161 , 
        \tx_fifo/n160 , \tx_fifo/n159 , \tx_fifo/n158 , \tx_fifo/n157 , 
        \tx_fifo/n156 , \tx_fifo/n155 , \data_to_tx_packet_len_reg[1] , 
        \data_to_tx_packet_len_reg[2] , \data_to_tx_packet_len_reg[3] , 
        \data_to_tx_packet_len_reg[4] , \data_to_tx_packet_len_reg[5] , 
        \data_to_tx_packet_len_reg[6] , \data_to_tx_packet_len_reg[7] , 
        \tx_fifo/n143 , \tx_fifo/n142 , \tx_fifo/n141 , \tx_fifo/n140 , 
        \tx_fifo/n139 , \tx_fifo/n138 , \tx_fifo/n137 , \rx_fifo/n153 , 
        ceg_net322, \rx_fifo/n162 , ceg_net340, \data_to_rx_packet_len_reg[0] , 
        rx_en_rx_packet_len, rx_en_rx_packet, \rx_fifo/n144 , ceg_net498, 
        \rx_fifo/n152 , \rx_fifo/n151 , \rx_fifo/n150 , \rx_fifo/n149 , 
        \rx_fifo/n148 , \rx_fifo/n147 , \rx_fifo/n146 , \rx_fifo/n161 , 
        \rx_fifo/n160 , \rx_fifo/n159 , \rx_fifo/n158 , \rx_fifo/n157 , 
        \rx_fifo/n156 , \rx_fifo/n155 , \data_to_rx_packet_len_reg[1] , 
        \data_to_rx_packet_len_reg[2] , \data_to_rx_packet_len_reg[3] , 
        \data_to_rx_packet_len_reg[4] , \data_to_rx_packet_len_reg[5] , 
        \data_to_rx_packet_len_reg[6] , \data_to_rx_packet_len_reg[7] , 
        \rx_fifo/n143 , \rx_fifo/n142 , \rx_fifo/n141 , \rx_fifo/n140 , 
        \rx_fifo/n139 , \rx_fifo/n138 , \rx_fifo/n137 , \i14/n128 , 
        \i14/n127 , \i14/n126 , \i14/n125 , \i14/n124 , \i14/n123 , 
        \i14/n122 , \i14/n121 , \i14/n120 , \i14/n119 , \i14/n118 , 
        \i14/n117 , \i14/n116 , \i14/n115 , \i14/n114 , \i14/n113 , 
        \i14/n112 , \i14/n111 , \i14/n110 , \i14/n109 , \i14/n108 , 
        \i14/n107 , \i14/n106 , \i14/n105 , \i14/n104 , \i14/n103 , 
        \i14/n102 , \i14/n101 , \i14/n100 , \i14/n99 , \i14/n98 , 
        \i14/n97 , \i14/n96 , \i14/n95 , \i14/n94 , \i14/n93 , \i14/n92 , 
        \i14/n91 , \i14/n90 , \i14/n89 , \i14/n88 , \i14/n87 , \i14/n86 , 
        \i14/n85 , \i14/n84 , \i14/n83 , \i14/n82 , \i14/n81 , \i14/n80 , 
        \i14/n79 , \i14/n78 , \i14/n77 , \i14/n76 , \i14/n75 , \i14/n74 , 
        \i14/n73 , \i14/n72 , \i14/n71 , \i14/n70 , \i14/n69 , \i14/n68 , 
        \i14/n67 , \i14/n66 , \i14/n65 , \i14/n64 , \i14/n63 , \i14/n62 , 
        \i14/n61 , \i14/n60 , \i14/n59 , \i14/n58 , \i14/n57 , \i14/n56 , 
        \i14/n55 , \i14/n54 , \i14/n53 , \i14/n52 , \i14/n51 , \i14/n50 , 
        \i14/n49 , \i14/n48 , \i14/n47 , \i14/n46 , \i14/n45 , \i14/n44 , 
        \i14/n43 , \i14/n42 , \i14/n41 , \i14/n40 , \i14/n39 , \i14/n38 , 
        \i14/n37 , \i14/n36 , \i14/n35 , \i14/n34 , \i14/n33 , \i14/n32 , 
        \i14/n31 , \i14/n30 , \i14/n29 , \i14/n28 , \i14/n27 , \i14/n26 , 
        \i14/n25 , \i14/n24 , \i14/n23 , \i14/n22 , \i14/n21 , \i14/n20 , 
        \i14/n19 , \i14/n18 , \i14/n17 , \i14/n16 , \i14/n15 , \i14/n14 , 
        \i14/n13 , \i14/n12 , \i14/n11 , \i14/n10 , \i14/n9 , \i14/n8 , 
        \i14/n7 , \i14/n6 , \i14/n5 , \data_to_tx_packet_reg[0] , \i15/n132 , 
        \data_to_tx_packet_reg[1] , \data_to_tx_packet_reg[2] , \data_to_tx_packet_reg[3] , 
        \data_to_tx_packet_reg[4] , \data_to_tx_packet_reg[5] , \data_to_tx_packet_reg[6] , 
        \data_to_tx_packet_reg[7] , \i15/n131 , \i15/n130 , \i15/n129 , 
        \i15/n128 , \i15/n127 , \i15/n126 , \i15/n125 , \i15/n124 , 
        \i15/n123 , \i15/n122 , \i15/n121 , \i15/n120 , \i15/n119 , 
        \i15/n118 , \i15/n117 , \i15/n116 , \i15/n115 , \i15/n114 , 
        \i15/n113 , \i15/n112 , \i15/n111 , \i15/n110 , \i15/n109 , 
        \i15/n108 , \i15/n107 , \i15/n106 , \i15/n105 , \i15/n104 , 
        \i15/n103 , \i15/n102 , \i15/n101 , \i15/n100 , \i15/n99 , 
        \i15/n98 , \i15/n97 , \i15/n96 , \i15/n95 , \i15/n94 , \i15/n93 , 
        \i15/n92 , \i15/n91 , \i15/n90 , \i15/n89 , \i15/n88 , \i15/n87 , 
        \i15/n86 , \i15/n85 , \i15/n84 , \i15/n83 , \i15/n82 , \i15/n81 , 
        \i15/n80 , \i15/n79 , \i15/n78 , \i15/n77 , \i15/n76 , \i15/n75 , 
        \i15/n74 , \i15/n73 , \i15/n72 , \i15/n71 , \i15/n70 , \i15/n69 , 
        \i15/n68 , \i15/n67 , \i15/n66 , \i15/n65 , \i15/n64 , \i15/n63 , 
        \i15/n62 , \i15/n61 , \i15/n60 , \i15/n59 , \i15/n58 , \i15/n57 , 
        \i15/n56 , \i15/n55 , \i15/n54 , \i15/n53 , \i15/n52 , \i15/n51 , 
        \i15/n50 , \i15/n49 , \i15/n48 , \i15/n47 , \i15/n46 , \i15/n45 , 
        \i15/n44 , \i15/n43 , \i15/n42 , \i15/n41 , \i15/n40 , \i15/n39 , 
        \i15/n38 , \i15/n37 , \i15/n36 , \i15/n35 , \i15/n34 , \i15/n33 , 
        \i15/n32 , \i15/n31 , \i15/n30 , \i15/n29 , \i15/n28 , \i15/n27 , 
        \i15/n26 , \i15/n25 , \i15/n24 , \i15/n23 , \i15/n22 , \i15/n21 , 
        \i15/n20 , \i15/n19 , \i15/n18 , \i15/n17 , \i15/n16 , \i15/n15 , 
        \i15/n14 , \i15/n13 , \i15/n12 , \i15/n11 , \i15/n10 , \i15/n9 , 
        \i15/n8 , \i15/n7 , \i15/n6 , \i15/n5 , \data_to_rx_packet_reg[0] , 
        \i16/n132 , \data_to_rx_packet_reg[1] , \data_to_rx_packet_reg[2] , 
        \data_to_rx_packet_reg[3] , \data_to_rx_packet_reg[4] , \data_to_rx_packet_reg[5] , 
        \data_to_rx_packet_reg[6] , \data_to_rx_packet_reg[7] , \i16/n131 , 
        \i16/n130 , \i16/n129 , \i16/n128 , \i16/n127 , \i16/n126 , 
        \i16/n125 , \i16/n124 , \i16/n123 , \i16/n122 , \i16/n121 , 
        \i16/n120 , \i16/n119 , \i16/n118 , \i16/n117 , \i16/n116 , 
        \i16/n115 , \i16/n114 , \i16/n113 , \i16/n112 , \i16/n111 , 
        \i16/n110 , \i16/n109 , \i16/n108 , \i16/n107 , \i16/n106 , 
        \i16/n105 , \i16/n104 , \i16/n103 , \i16/n102 , \i16/n101 , 
        \i16/n100 , \i16/n99 , \i16/n98 , \i16/n97 , \i16/n96 , \i16/n95 , 
        \i16/n94 , \i16/n93 , \i16/n92 , \i16/n91 , \i16/n90 , \i16/n89 , 
        \i16/n88 , \i16/n87 , \i16/n86 , \i16/n85 , \i16/n84 , \i16/n83 , 
        \i16/n82 , \i16/n81 , \i16/n80 , \i16/n79 , \i16/n78 , \i16/n77 , 
        \i16/n76 , \i16/n75 , \i16/n74 , \i16/n73 , \i16/n72 , \i16/n71 , 
        \i16/n70 , \i16/n69 , \i16/n68 , \i16/n67 , \i16/n66 , \i16/n65 , 
        \i16/n64 , \i16/n63 , \i16/n62 , \i16/n61 , \i16/n60 , \i16/n59 , 
        \i16/n58 , \i16/n57 , \i16/n56 , \i16/n55 , \i16/n54 , \i16/n53 , 
        \i16/n52 , \i16/n51 , \i16/n50 , \i16/n49 , \i16/n48 , \i16/n47 , 
        \i16/n46 , \i16/n45 , \i16/n44 , \i16/n43 , \i16/n42 , \i16/n41 , 
        \i16/n40 , \i16/n39 , \i16/n38 , \i16/n37 , \i16/n36 , \i16/n35 , 
        \i16/n34 , \i16/n33 , \i16/n32 , \i16/n31 , \i16/n30 , \i16/n29 , 
        \i16/n28 , \i16/n27 , \i16/n26 , \i16/n25 , \i16/n24 , \i16/n23 , 
        \i16/n22 , \i16/n21 , \i16/n20 , \i16/n19 , \i16/n18 , \i16/n17 , 
        \i16/n16 , n4152, \i16/n15 , n4161, \i16/n14 , \i16/n13 , 
        n4167, \i16/n12 , \i16/n11 , \i16/n10 , \i16/n9 , \i16/n8 , 
        \i16/n7 , \i16/n6 , \i16/n5 , \pll_clk~O , \tx_slowclk~O , 
        n7059, n7058, n7057, n7056, n7055, n4235, n4236, n4237, 
        n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, 
        n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, 
        n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, 
        n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, 
        n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, 
        n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, 
        n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, 
        n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, 
        n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, 
        n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, 
        n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, 
        n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, 
        n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, 
        n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, 
        n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, 
        n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, 
        n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, 
        n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, 
        n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, 
        n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, 
        n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, 
        n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, 
        n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, 
        n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, 
        n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, 
        n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, 
        n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, 
        n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, 
        n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, 
        n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, 
        n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, 
        n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, 
        n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, 
        n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, 
        n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, 
        n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, 
        n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, 
        n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, 
        n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, 
        n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, 
        n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, 
        n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, 
        n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, 
        n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, 
        n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, 
        n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, 
        n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, 
        n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, 
        n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, 
        n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, 
        n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, 
        n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, 
        n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, 
        n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, 
        n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, 
        n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, 
        n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, 
        n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, 
        n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, 
        n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, 
        n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, 
        n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, 
        n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, 
        n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, 
        n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, 
        n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, 
        n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, 
        n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, 
        n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, 
        n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, 
        n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, 
        n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, 
        n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, 
        n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, 
        n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, 
        n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, 
        n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, 
        n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, 
        n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, 
        n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, 
        n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, 
        n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, 
        n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, 
        n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, 
        n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, 
        n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, 
        n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, 
        n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, 
        n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, 
        n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, 
        n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, 
        n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, 
        n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, 
        n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, 
        n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, 
        n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, 
        n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, 
        n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, 
        n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, 
        n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, 
        n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, 
        n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, 
        n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, 
        n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, 
        n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, 
        n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, 
        n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, 
        n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, 
        n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, 
        n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, 
        n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, 
        n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, 
        n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, 
        n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, 
        n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, 
        n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, 
        n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, 
        n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, 
        n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, 
        n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, 
        n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, 
        n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, 
        n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, 
        n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, 
        n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, 
        n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, 
        n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, 
        n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, 
        n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, 
        n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, 
        n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, 
        n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, 
        n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, 
        n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, 
        n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, 
        n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, 
        n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, 
        n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, 
        n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, 
        n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, 
        n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, 
        n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, 
        n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, 
        n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, 
        n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, 
        n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, 
        n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, 
        n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, 
        n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, 
        n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, 
        n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, 
        n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, 
        n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, 
        n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, 
        n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, 
        n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, 
        n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, 
        n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, 
        n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, 
        n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, 
        n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, 
        n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, 
        n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, 
        n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, 
        n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, 
        n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, 
        n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, 
        n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, 
        n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, 
        n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, 
        n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, 
        n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, 
        n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, 
        n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, 
        n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, 
        n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, 
        n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, 
        n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, 
        n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, 
        n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, 
        n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, 
        n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, 
        n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, 
        n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, 
        n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, 
        n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, 
        n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, 
        n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, 
        n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, 
        n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, 
        n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, 
        n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, 
        n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, 
        n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, 
        n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, 
        n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, 
        n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, 
        n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, 
        n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, 
        n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, 
        n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, 
        n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, 
        n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, 
        n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, 
        n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, 
        n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, 
        n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, 
        n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, 
        n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, 
        n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, 
        n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, 
        n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, 
        n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, 
        n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, 
        n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, 
        n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, 
        n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, 
        n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, 
        n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, 
        n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, 
        n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, 
        n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, 
        n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, 
        n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, 
        n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, 
        n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, 
        n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, 
        n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, 
        n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, 
        n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, 
        n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, 
        n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, 
        n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, 
        n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, 
        n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, 
        n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, 
        n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, 
        n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, 
        n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, 
        n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, 
        n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, 
        n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, 
        n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, 
        n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, 
        n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, 
        n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, 
        n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, 
        n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, 
        n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, 
        n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, 
        n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, 
        n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, 
        n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, 
        n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, 
        n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, 
        n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, 
        n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, 
        n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, 
        n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, 
        n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, 
        n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, 
        n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, 
        n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, 
        n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, 
        n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, 
        n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, 
        n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, 
        n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, 
        n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, 
        n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, 
        n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, 
        n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, 
        n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, 
        n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, 
        n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, 
        n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, 
        n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, 
        n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, 
        n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, 
        n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, 
        n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, 
        n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, 
        n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, 
        n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, 
        n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, 
        n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, 
        n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, 
        n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, 
        n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, 
        n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, 
        n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, 
        n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, 
        n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, 
        n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, 
        n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, 
        n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, 
        n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, 
        n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, 
        n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, 
        n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, 
        n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, 
        n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, 
        n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, 
        n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, 
        n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, 
        n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, 
        n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, 
        n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, 
        n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, 
        n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, 
        n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, 
        n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, 
        n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, 
        n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, 
        n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, 
        n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, 
        n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, 
        n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, 
        n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, 
        n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, 
        n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, 
        n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, 
        n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, 
        n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, 
        n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, 
        n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, 
        n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, 
        n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, 
        n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, 
        n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, 
        n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, 
        n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, 
        n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, 
        n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, 
        n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, 
        n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, 
        n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, 
        n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, 
        n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, 
        n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, 
        n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, 
        n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, 
        n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, 
        n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, 
        n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, 
        n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, 
        n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, 
        n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, 
        n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, 
        n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, 
        n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, 
        n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, 
        n7054;
    
    EFX_LUT4 \tx_dac_fsm_inst/i116  (.I0(n3561), .I1(n113), .I2(n3562), 
            .O(n113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/i116 .LUTMASK = 16'hacac;
    EFX_FF \reg_addr[4]~FF  (.D(\spi_slave_inst/n94 ), .CE(ceg_net49), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\reg_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(114)
    defparam \reg_addr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \reg_addr[4]~FF .CE_POLARITY = 1'b0;
    defparam \reg_addr[4]~FF .SR_POLARITY = 1'b0;
    defparam \reg_addr[4]~FF .D_POLARITY = 1'b1;
    defparam \reg_addr[4]~FF .SR_SYNC = 1'b0;
    defparam \reg_addr[4]~FF .SR_VALUE = 1'b0;
    defparam \reg_addr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \reg_addr[3]~FF  (.D(\spi_slave_inst/n95 ), .CE(ceg_net49), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\reg_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(114)
    defparam \reg_addr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \reg_addr[3]~FF .CE_POLARITY = 1'b0;
    defparam \reg_addr[3]~FF .SR_POLARITY = 1'b0;
    defparam \reg_addr[3]~FF .D_POLARITY = 1'b1;
    defparam \reg_addr[3]~FF .SR_SYNC = 1'b0;
    defparam \reg_addr[3]~FF .SR_VALUE = 1'b0;
    defparam \reg_addr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/bitcnt[2]~FF  (.D(\spi_slave_inst/n56 ), .CE(ceg_net40), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/bitcnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/bitcnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[2]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[2]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/bitcnt[2]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/bitcnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/bitcnt[1]~FF  (.D(\spi_slave_inst/n57 ), .CE(ceg_net40), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/bitcnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/bitcnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[1]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[1]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/bitcnt[1]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/bitcnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_tx_en[1]~FF  (.D(\spi_slave_inst/sync_tx_en[0] ), 
           .CE(1'b1), .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/sync_tx_en[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_tx_en[1]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_tx_en[1]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_tx_en[1]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_tx_en[1]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_tx_en[1]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_tx_en[1]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/sync_tx_en[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \reg_addr[2]~FF  (.D(\spi_slave_inst/n96 ), .CE(ceg_net49), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\reg_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(114)
    defparam \reg_addr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \reg_addr[2]~FF .CE_POLARITY = 1'b0;
    defparam \reg_addr[2]~FF .SR_POLARITY = 1'b0;
    defparam \reg_addr[2]~FF .D_POLARITY = 1'b1;
    defparam \reg_addr[2]~FF .SR_SYNC = 1'b0;
    defparam \reg_addr[2]~FF .SR_VALUE = 1'b0;
    defparam \reg_addr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \reg_addr[1]~FF  (.D(\spi_slave_inst/n97 ), .CE(ceg_net49), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\reg_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(114)
    defparam \reg_addr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \reg_addr[1]~FF .CE_POLARITY = 1'b0;
    defparam \reg_addr[1]~FF .SR_POLARITY = 1'b0;
    defparam \reg_addr[1]~FF .D_POLARITY = 1'b1;
    defparam \reg_addr[1]~FF .SR_SYNC = 1'b0;
    defparam \reg_addr[1]~FF .SR_VALUE = 1'b0;
    defparam \reg_addr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_tx_en[0]_2~FF  (.D(tx_en), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\spi_slave_inst/sync_tx_en[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_tx_en[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_tx_en[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_tx_en[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_tx_en[0]_2~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_tx_en[0]_2~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_tx_en[0]_2~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/sync_tx_en[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/bitcnt[0]~FF  (.D(\spi_slave_inst/n58 ), .CE(ceg_net40), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/bitcnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/bitcnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[0]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[0]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/bitcnt[0]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/bitcnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_mosi[1]~FF  (.D(\spi_slave_inst/sync_mosi[0] ), 
           .CE(1'b1), .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/sync_mosi[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_mosi[1]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_mosi[1]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_mosi[1]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_mosi[1]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_mosi[1]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_mosi[1]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/sync_mosi[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rw_out~FF  (.D(\spi_slave_inst/n73 ), .CE(ceg_net23), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(rw_out)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(103)
    defparam \rw_out~FF .CLK_POLARITY = 1'b1;
    defparam \rw_out~FF .CE_POLARITY = 1'b0;
    defparam \rw_out~FF .SR_POLARITY = 1'b0;
    defparam \rw_out~FF .D_POLARITY = 1'b1;
    defparam \rw_out~FF .SR_SYNC = 1'b0;
    defparam \rw_out~FF .SR_VALUE = 1'b0;
    defparam \rw_out~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \reg_addr[0]~FF  (.D(\spi_slave_inst/n98 ), .CE(ceg_net49), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\reg_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(114)
    defparam \reg_addr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \reg_addr[0]~FF .CE_POLARITY = 1'b0;
    defparam \reg_addr[0]~FF .SR_POLARITY = 1'b0;
    defparam \reg_addr[0]~FF .D_POLARITY = 1'b1;
    defparam \reg_addr[0]~FF .SR_SYNC = 1'b0;
    defparam \reg_addr[0]~FF .SR_VALUE = 1'b0;
    defparam \reg_addr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[0]~FF  (.D(\spi_slave_inst/n139 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[0]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[0]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[0]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[0]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[0]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[0]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[0]~FF  (.D(\spi_slave_inst/n98 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[0]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[0]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[0]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[0]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[0]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[0]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \addr_dv~FF  (.D(\spi_slave_inst/n68 ), .CE(ceg_net34), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(addr_dv)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(155)
    defparam \addr_dv~FF .CLK_POLARITY = 1'b1;
    defparam \addr_dv~FF .CE_POLARITY = 1'b0;
    defparam \addr_dv~FF .SR_POLARITY = 1'b0;
    defparam \addr_dv~FF .D_POLARITY = 1'b0;
    defparam \addr_dv~FF .SR_SYNC = 1'b0;
    defparam \addr_dv~FF .SR_VALUE = 1'b0;
    defparam \addr_dv~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rxdv~FF  (.D(\spi_slave_inst/n68 ), .CE(ceg_net37), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(rxdv)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(165)
    defparam \rxdv~FF .CLK_POLARITY = 1'b1;
    defparam \rxdv~FF .CE_POLARITY = 1'b0;
    defparam \rxdv~FF .SR_POLARITY = 1'b0;
    defparam \rxdv~FF .D_POLARITY = 1'b0;
    defparam \rxdv~FF .SR_SYNC = 1'b0;
    defparam \rxdv~FF .SR_VALUE = 1'b0;
    defparam \rxdv~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_sclk[0]~FF  (.D(SCLK), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\spi_slave_inst/sync_sclk[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_sclk[0]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[0]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[0]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_sclk[0]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[0]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_sclk[0]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/sync_sclk[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/bitcnt[4]~FF  (.D(\spi_slave_inst/n54 ), .CE(ceg_net40), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/bitcnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/bitcnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[4]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[4]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/bitcnt[4]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/bitcnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \reg_addr[5]~FF  (.D(\spi_slave_inst/n93 ), .CE(ceg_net49), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\reg_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(114)
    defparam \reg_addr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \reg_addr[5]~FF .CE_POLARITY = 1'b0;
    defparam \reg_addr[5]~FF .SR_POLARITY = 1'b0;
    defparam \reg_addr[5]~FF .D_POLARITY = 1'b1;
    defparam \reg_addr[5]~FF .SR_SYNC = 1'b0;
    defparam \reg_addr[5]~FF .SR_VALUE = 1'b0;
    defparam \reg_addr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/bitcnt[3]~FF  (.D(\spi_slave_inst/n55 ), .CE(ceg_net40), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/bitcnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/bitcnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/bitcnt[3]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/bitcnt[3]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/bitcnt[3]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/bitcnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_mosi[0]_2~FF  (.D(MOSI), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\spi_slave_inst/sync_mosi[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_mosi[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_mosi[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_mosi[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_mosi[0]_2~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_mosi[0]_2~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_mosi[0]_2~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/sync_mosi[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_ss[0]~FF  (.D(SSB), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\spi_slave_inst/sync_ss[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_ss[0]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[0]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[0]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_ss[0]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[0]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_ss[0]~FF .SR_VALUE = 1'b1;
    defparam \spi_slave_inst/sync_ss[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \reg_addr[6]~FF  (.D(\spi_slave_inst/n92 ), .CE(ceg_net49), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\reg_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(114)
    defparam \reg_addr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \reg_addr[6]~FF .CE_POLARITY = 1'b0;
    defparam \reg_addr[6]~FF .SR_POLARITY = 1'b0;
    defparam \reg_addr[6]~FF .D_POLARITY = 1'b1;
    defparam \reg_addr[6]~FF .SR_SYNC = 1'b0;
    defparam \reg_addr[6]~FF .SR_VALUE = 1'b0;
    defparam \reg_addr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[1]~FF  (.D(\spi_slave_inst/n138 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[1]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[1]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[1]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[1]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[1]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[2]~FF  (.D(\spi_slave_inst/n137 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[2]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[2]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[2]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[2]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[2]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[2]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[3]~FF  (.D(\spi_slave_inst/n136 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[3]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[3]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[3]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[3]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[3]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[3]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[4]~FF  (.D(\spi_slave_inst/n135 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[4]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[4]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[4]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[4]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[4]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[4]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[5]~FF  (.D(\spi_slave_inst/n134 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[5]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[5]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[5]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[5]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[5]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[5]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[6]~FF  (.D(\spi_slave_inst/n133 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[6]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[6]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[6]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[6]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[6]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[6]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/d_o[7]~FF  (.D(\spi_slave_inst/n132 ), .CE(ceg_net77), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/d_o[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(132)
    defparam \spi_slave_inst/d_o[7]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[7]~FF .CE_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[7]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/d_o[7]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/d_o[7]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/d_o[7]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/d_o[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[1]~FF  (.D(\spi_slave_inst/n173 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[1]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[1]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[1]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[1]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[1]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[1]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[2]~FF  (.D(\spi_slave_inst/n172 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[2]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[2]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[2]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[2]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[2]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[2]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[3]~FF  (.D(\spi_slave_inst/n171 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[3]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[3]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[3]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[3]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[3]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[3]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[4]~FF  (.D(\spi_slave_inst/n170 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[4]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[4]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[4]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[4]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[4]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[4]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[5]~FF  (.D(\spi_slave_inst/n169 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[5]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[5]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[5]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[5]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[5]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[5]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[6]~FF  (.D(\spi_slave_inst/n168 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[6]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[6]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[6]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[6]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[6]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[6]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_d[7]~FF  (.D(\spi_slave_inst/n167 ), .CE(ceg_net98), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_d[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(143)
    defparam \rx_d[7]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_d[7]~FF .CE_POLARITY = 1'b0;
    defparam \rx_d[7]~FF .SR_POLARITY = 1'b0;
    defparam \rx_d[7]~FF .D_POLARITY = 1'b1;
    defparam \rx_d[7]~FF .SR_SYNC = 1'b0;
    defparam \rx_d[7]~FF .SR_VALUE = 1'b0;
    defparam \rx_d[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_sclk[1]~FF  (.D(\spi_slave_inst/sync_sclk[0] ), 
           .CE(1'b1), .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/sync_sclk[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_sclk[1]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[1]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[1]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_sclk[1]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[1]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_sclk[1]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/sync_sclk[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_sclk[2]~FF  (.D(\spi_slave_inst/sync_sclk[1] ), 
           .CE(1'b1), .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/sync_sclk[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_sclk[2]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[2]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[2]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_sclk[2]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_sclk[2]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_sclk[2]~FF .SR_VALUE = 1'b0;
    defparam \spi_slave_inst/sync_sclk[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_ss[1]~FF  (.D(\spi_slave_inst/sync_ss[0] ), 
           .CE(1'b1), .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/sync_ss[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_ss[1]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[1]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[1]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_ss[1]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[1]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_ss[1]~FF .SR_VALUE = 1'b1;
    defparam \spi_slave_inst/sync_ss[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \spi_slave_inst/sync_ss[2]~FF  (.D(\spi_slave_inst/sync_ss[1] ), 
           .CE(1'b1), .CLK(\pll_clk~O ), .SR(reset_n), .Q(\spi_slave_inst/sync_ss[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(62)
    defparam \spi_slave_inst/sync_ss[2]~FF .CLK_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[2]~FF .CE_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[2]~FF .SR_POLARITY = 1'b0;
    defparam \spi_slave_inst/sync_ss[2]~FF .D_POLARITY = 1'b1;
    defparam \spi_slave_inst/sync_ss[2]~FF .SR_SYNC = 1'b0;
    defparam \spi_slave_inst/sync_ss[2]~FF .SR_VALUE = 1'b1;
    defparam \spi_slave_inst/sync_ss[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[7]~FF  (.D(\led_inst/n41 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[7]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[7]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[7]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[7]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[7]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[7]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[6]~FF  (.D(\led_inst/n42 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[6]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[6]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[6]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[6]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[6]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[6]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[5]~FF  (.D(\led_inst/n43 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[5]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[5]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[5]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[5]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[5]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[5]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[4]~FF  (.D(\led_inst/n44 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[4]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[4]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[4]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[4]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[4]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[4]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[3]~FF  (.D(\led_inst/n45 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[3]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[3]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[3]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[3]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[3]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[3]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[0]~FF  (.D(\led_inst/n48 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[0]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[0]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[0]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[0]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[0]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[0]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[2]~FF  (.D(\led_inst/n46 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[2]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[2]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[2]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[2]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[2]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[2]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_from_led[1]~FF  (.D(\led_inst/n47 ), .CE(1'b0), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\data_from_led[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(58)
    defparam \data_from_led[1]~FF .CLK_POLARITY = 1'b1;
    defparam \data_from_led[1]~FF .CE_POLARITY = 1'b0;
    defparam \data_from_led[1]~FF .SR_POLARITY = 1'b0;
    defparam \data_from_led[1]~FF .D_POLARITY = 1'b1;
    defparam \data_from_led[1]~FF .SR_SYNC = 1'b0;
    defparam \data_from_led[1]~FF .SR_VALUE = 1'b0;
    defparam \data_from_led[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[0]~FF  (.D(\led_inst/n142 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[0]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[0]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[0]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[0]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[0]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[0]~FF  (.D(\data_to_led[0] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[0]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[0]~FF .SR_VALUE = 1'b1;
    defparam \led_inst/ctr_cfg_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led0~FF  (.D(led0), .CE(\led_inst/LessThan_21/n48 ), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(led0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led0~FF .CLK_POLARITY = 1'b1;
    defparam \led0~FF .CE_POLARITY = 1'b1;
    defparam \led0~FF .SR_POLARITY = 1'b0;
    defparam \led0~FF .D_POLARITY = 1'b0;
    defparam \led0~FF .SR_SYNC = 1'b0;
    defparam \led0~FF .SR_VALUE = 1'b0;
    defparam \led0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led1~FF  (.D(led0), .CE(\led_inst/LessThan_21/n48 ), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(led1)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led1~FF .CLK_POLARITY = 1'b1;
    defparam \led1~FF .CE_POLARITY = 1'b1;
    defparam \led1~FF .SR_POLARITY = 1'b0;
    defparam \led1~FF .D_POLARITY = 1'b1;
    defparam \led1~FF .SR_SYNC = 1'b0;
    defparam \led1~FF .SR_VALUE = 1'b1;
    defparam \led1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[1]~FF  (.D(\led_inst/n141 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[1]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[1]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[1]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[1]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[2]~FF  (.D(\led_inst/n140 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[2]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[2]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[2]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[2]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[3]~FF  (.D(\led_inst/n139 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[3]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[3]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[3]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[3]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[4]~FF  (.D(\led_inst/n138 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[4]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[4]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[4]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[4]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[5]~FF  (.D(\led_inst/n137 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[5]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[5]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[5]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[5]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[6]~FF  (.D(\led_inst/n136 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[6]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[6]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[6]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[6]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[6]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[7]~FF  (.D(\led_inst/n135 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[7]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[7]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[7]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[7]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[7]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[8]~FF  (.D(\led_inst/n134 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[8]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[8]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[8]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[8]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[8]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[9]~FF  (.D(\led_inst/n133 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[9]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[9]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[9]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[9]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[9]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[10]~FF  (.D(\led_inst/n132 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[10]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[10]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[10]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[10]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[10]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[11]~FF  (.D(\led_inst/n131 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[11]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[11]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[11]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[11]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[11]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[12]~FF  (.D(\led_inst/n130 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[12]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[12]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[12]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[12]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[12]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[13]~FF  (.D(\led_inst/n129 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[13]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[13]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[13]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[13]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[13]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[14]~FF  (.D(\led_inst/n128 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[14]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[14]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[14]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[14]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[14]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[15]~FF  (.D(\led_inst/n127 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[15]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[15]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[15]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[15]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[15]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[16]~FF  (.D(\led_inst/n126 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[16]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[16]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[16]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[16]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[16]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[16]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[17]~FF  (.D(\led_inst/n125 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[17]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[17]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[17]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[17]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[17]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[17]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[18]~FF  (.D(\led_inst/n124 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[18]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[18]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[18]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[18]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[18]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[18]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[19]~FF  (.D(\led_inst/n123 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[19]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[19]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[19]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[19]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[19]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[19]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[20]~FF  (.D(\led_inst/n122 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[20]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[20]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[20]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[20]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[20]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[20]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[21]~FF  (.D(\led_inst/n121 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[21]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[21]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[21]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[21]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[21]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[21]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[22]~FF  (.D(\led_inst/n120 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[22]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[22]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[22]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[22]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[22]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[22]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/counter[23]~FF  (.D(\led_inst/n119 ), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\led_inst/counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(79)
    defparam \led_inst/counter[23]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/counter[23]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/counter[23]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/counter[23]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/counter[23]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/counter[23]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/counter[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[1]~FF  (.D(\data_to_led[1] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[1]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/ctr_cfg_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[2]~FF  (.D(\data_to_led[2] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[2]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[2]~FF .SR_VALUE = 1'b1;
    defparam \led_inst/ctr_cfg_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[3]~FF  (.D(\data_to_led[3] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[3]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[3]~FF .SR_VALUE = 1'b1;
    defparam \led_inst/ctr_cfg_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[4]~FF  (.D(\data_to_led[4] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[4]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[4]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[4]~FF .SR_VALUE = 1'b1;
    defparam \led_inst/ctr_cfg_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[5]~FF  (.D(\data_to_led[5] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[5]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[5]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/ctr_cfg_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[6]~FF  (.D(\data_to_led[6] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[6]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[6]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[6]~FF .SR_VALUE = 1'b1;
    defparam \led_inst/ctr_cfg_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_inst/ctr_cfg_reg[7]~FF  (.D(\data_to_led[7] ), .CE(rx_en_led), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\led_inst/ctr_cfg_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(46)
    defparam \led_inst/ctr_cfg_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[7]~FF .CE_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[7]~FF .SR_POLARITY = 1'b0;
    defparam \led_inst/ctr_cfg_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \led_inst/ctr_cfg_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \led_inst/ctr_cfg_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \led_inst/ctr_cfg_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[0]~FF  (.D(\data_to_gpo[0] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[0]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[1]~FF  (.D(\data_to_gpo[1] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[1]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[2]~FF  (.D(\data_to_gpo[2] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[2]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[3]~FF  (.D(\data_to_gpo[3] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[3]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[4]~FF  (.D(\data_to_gpo[4] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[4]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[4]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[5]~FF  (.D(\data_to_gpo[5] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[5]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[5]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[6]~FF  (.D(\data_to_gpo[6] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[6]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[6]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \gpo_inst/gp_config_reg[7]~FF  (.D(\data_to_gpo[7] ), .CE(rx_en_gpo), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\gpo_inst/gp_config_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\gpo.sv(21)
    defparam \gpo_inst/gp_config_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[7]~FF .CE_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[7]~FF .SR_POLARITY = 1'b0;
    defparam \gpo_inst/gp_config_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \gpo_inst/gp_config_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \gpo_inst/gp_config_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \gpo_inst/gp_config_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[3][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[3][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[3][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[3][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[3][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[3][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[3][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[3][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[3][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[3][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[3][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[3][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[3][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[3][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[3][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[2][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[2][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[2][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[2][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[2][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_ctr[0]~FF  (.D(\tx_dac_fsm_inst/n68 ), .CE(\tx_dac_fsm_inst/n42 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_ctr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_ctr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_pos[0]~FF  (.D(\tx_dac_fsm_inst/sym_pos[0] ), 
           .CE(\tx_dac_fsm_inst/n344 ), .CLK(\tx_slowclk~O ), .SR(reset_n), 
           .Q(\tx_dac_fsm_inst/sym_pos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_pos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[0]~FF .D_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/state_reg[0]~FF  (.D(n109), .CE(1'b1), .CLK(\tx_slowclk~O ), 
           .SR(reset_n), .Q(\tx_dac_fsm_inst/state_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(113)
    defparam \tx_dac_fsm_inst/state_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_ctr[1]~FF  (.D(\tx_dac_fsm_inst/n67 ), .CE(\tx_dac_fsm_inst/n42 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_ctr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_ctr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[1]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_ctr[2]~FF  (.D(\tx_dac_fsm_inst/n66 ), .CE(\tx_dac_fsm_inst/n42 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_ctr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_ctr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[2]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[2]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[2]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[2]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[2]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_ctr[3]~FF  (.D(\tx_dac_fsm_inst/n65 ), .CE(\tx_dac_fsm_inst/n42 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_ctr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_ctr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[3]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[3]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[3]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[3]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[3]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[2][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[2][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[2][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[2][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[2][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/zctr[0]~FF  (.D(\tx_dac_fsm_inst/n258 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/zctr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(200)
    defparam \tx_dac_fsm_inst/zctr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_ctr[4]~FF  (.D(\tx_dac_fsm_inst/n64 ), .CE(\tx_dac_fsm_inst/n42 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_ctr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_ctr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[4]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[4]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[4]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_ctr[4]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[4]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_ctr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dctr[0]~FF  (.D(\tx_dac_fsm_inst/n284 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/dctr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(211)
    defparam \tx_dac_fsm_inst/dctr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dac_config_reg[0]~FF  (.D(data_to_dac), .CE(rx_en_dac), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/dac_config_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(51)
    defparam \tx_dac_fsm_inst/dac_config_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dac_config_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dac_config_reg[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dac_config_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dac_config_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dac_config_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dac_config_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_pos[1]~FF  (.D(\~tx_dac_fsm_inst/n431 ), .CE(\tx_dac_fsm_inst/n344 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_pos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_pos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[1]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_pos[2]~FF  (.D(\~tx_dac_fsm_inst/n436 ), .CE(\tx_dac_fsm_inst/n344 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_pos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_pos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[2]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[2]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[2]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[2]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[2]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/sym_pos[3]~FF  (.D(\~tx_dac_fsm_inst/n441 ), .CE(\tx_dac_fsm_inst/n344 ), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/sym_pos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(103)
    defparam \tx_dac_fsm_inst/sym_pos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[3]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[3]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[3]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sym_pos[3]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[3]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/sym_pos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/state_reg[1]~FF  (.D(n133), .CE(1'b1), .CLK(\tx_slowclk~O ), 
           .SR(reset_n), .Q(\tx_dac_fsm_inst/state_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(113)
    defparam \tx_dac_fsm_inst/state_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/state_reg[2]~FF  (.D(n134), .CE(1'b1), .CLK(\tx_slowclk~O ), 
           .SR(reset_n), .Q(\tx_dac_fsm_inst/state_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(113)
    defparam \tx_dac_fsm_inst/state_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[2]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/state_reg[3]~FF  (.D(n135), .CE(1'b1), .CLK(\tx_slowclk~O ), 
           .SR(reset_n), .Q(\tx_dac_fsm_inst/state_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(113)
    defparam \tx_dac_fsm_inst/state_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[3]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/state_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/state_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/zctr[1]~FF  (.D(\tx_dac_fsm_inst/n257 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/zctr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(200)
    defparam \tx_dac_fsm_inst/zctr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[1]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/zctr[2]~FF  (.D(\tx_dac_fsm_inst/n256 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/zctr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(200)
    defparam \tx_dac_fsm_inst/zctr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[2]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[2]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[2]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[2]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[2]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/zctr[3]~FF  (.D(\tx_dac_fsm_inst/n255 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/zctr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(200)
    defparam \tx_dac_fsm_inst/zctr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[3]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[3]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[3]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[3]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[3]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/zctr[4]~FF  (.D(\tx_dac_fsm_inst/n254 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/zctr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(200)
    defparam \tx_dac_fsm_inst/zctr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[4]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[4]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[4]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[4]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[4]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/zctr[5]~FF  (.D(\tx_dac_fsm_inst/n253 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/zctr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(200)
    defparam \tx_dac_fsm_inst/zctr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[5]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[5]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[5]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/zctr[5]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[5]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/zctr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dctr[1]~FF  (.D(\tx_dac_fsm_inst/n283 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/dctr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(211)
    defparam \tx_dac_fsm_inst/dctr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[1]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dctr[2]~FF  (.D(\tx_dac_fsm_inst/n282 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/dctr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(211)
    defparam \tx_dac_fsm_inst/dctr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[2]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[2]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[2]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[2]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[2]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dctr[3]~FF  (.D(\tx_dac_fsm_inst/n281 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/dctr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(211)
    defparam \tx_dac_fsm_inst/dctr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[3]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[3]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[3]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[3]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[3]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dctr[4]~FF  (.D(\tx_dac_fsm_inst/n280 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/dctr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(211)
    defparam \tx_dac_fsm_inst/dctr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[4]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[4]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[4]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[4]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[4]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_dac_fsm_inst/dctr[5]~FF  (.D(\tx_dac_fsm_inst/n279 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(reset_n), .Q(\tx_dac_fsm_inst/dctr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(211)
    defparam \tx_dac_fsm_inst/dctr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[5]~FF .CE_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[5]~FF .SR_POLARITY = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[5]~FF .D_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/dctr[5]~FF .SR_SYNC = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[5]~FF .SR_VALUE = 1'b0;
    defparam \tx_dac_fsm_inst/dctr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[0]~FF  (.D(\fifo_inst/n153 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/wr_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[0]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[0]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[0]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[0]~FF  (.D(\fifo_inst/n162 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/rd_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[0]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[0]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[0]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[0]~FF  (.D(\data_to_fifo_length[0] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/length[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[0]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[0]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[0]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[0]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[0]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/sync_wr[0]~FF  (.D(rx_en_fifo), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\fifo_inst/sync_wr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/sync_wr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/sync_wr[0]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/sync_wr[0]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/sync_wr[0]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/sync_wr[0]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/sync_wr[0]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/sync_wr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/sync_rd[0]~FF  (.D(tx_en_fifo), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\fifo_inst/sync_rd[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/sync_rd[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/sync_rd[0]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/sync_rd[0]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/sync_rd[0]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/sync_rd[0]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/sync_rd[0]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/sync_rd[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[0]~FF  (.D(\fifo_inst/n144 ), .CE(ceg_net418), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/buff_head[0]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[0]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[0]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[0]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[0]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[0]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[1]~FF  (.D(\fifo_inst/n152 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/wr_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[1]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[1]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[1]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[2]~FF  (.D(\fifo_inst/n151 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/wr_index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[2]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[2]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[2]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[2]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[2]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[3]~FF  (.D(\fifo_inst/n150 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/wr_index[3]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[3]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[3]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[3]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[3]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[3]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[4]~FF  (.D(\fifo_inst/n149 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/wr_index[4]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[4]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[4]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[4]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[4]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[4]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[5]~FF  (.D(\fifo_inst/n148 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/wr_index[5]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[5]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[5]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[5]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[5]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[5]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[6]~FF  (.D(\fifo_inst/n147 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/wr_index[6]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[6]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[6]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[6]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[6]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[6]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/wr_index[7]~FF  (.D(\fifo_inst/n146 ), .CE(ceg_net146), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/wr_index[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/wr_index[7]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[7]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[7]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/wr_index[7]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/wr_index[7]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/wr_index[7]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/wr_index[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[1]~FF  (.D(\fifo_inst/n161 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/rd_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[1]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[1]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[1]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[2]~FF  (.D(\fifo_inst/n160 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/rd_index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[2]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[2]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[2]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[2]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[2]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[3]~FF  (.D(\fifo_inst/n159 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/rd_index[3]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[3]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[3]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[3]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[3]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[3]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[4]~FF  (.D(\fifo_inst/n158 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/rd_index[4]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[4]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[4]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[4]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[4]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[4]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[5]~FF  (.D(\fifo_inst/n157 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/rd_index[5]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[5]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[5]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[5]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[5]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[5]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[6]~FF  (.D(\fifo_inst/n156 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/rd_index[6]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[6]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[6]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[6]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[6]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[6]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/rd_index[7]~FF  (.D(\fifo_inst/n155 ), .CE(ceg_net164), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/rd_index[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/rd_index[7]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[7]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[7]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/rd_index[7]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/rd_index[7]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/rd_index[7]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/rd_index[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[1]~FF  (.D(\data_to_fifo_length[1] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/length[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[1]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[1]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[1]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[1]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[1]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[2]~FF  (.D(\data_to_fifo_length[2] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/length[2]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[2]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[2]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[2]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[2]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[2]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[3]~FF  (.D(\data_to_fifo_length[3] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/length[3]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[3]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[3]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[3]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[3]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[3]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[4]~FF  (.D(\data_to_fifo_length[4] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/length[4]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[4]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[4]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[4]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[4]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[4]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[5]~FF  (.D(\data_to_fifo_length[5] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/length[5]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[5]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[5]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[5]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[5]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[5]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[6]~FF  (.D(\data_to_fifo_length[6] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/length[6]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[6]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[6]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[6]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[6]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[6]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/length[7]~FF  (.D(\data_to_fifo_length[7] ), .CE(rx_en_fifo_length), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/length[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/length[7]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/length[7]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/length[7]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/length[7]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/length[7]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/length[7]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/length[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/sync_wr[1]~FF  (.D(\fifo_inst/sync_wr[0] ), .CE(1'b1), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/sync_wr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/sync_wr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/sync_wr[1]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/sync_wr[1]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/sync_wr[1]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/sync_wr[1]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/sync_wr[1]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/sync_wr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/sync_rd[1]~FF  (.D(\fifo_inst/sync_rd[0] ), .CE(1'b1), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/sync_rd[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/sync_rd[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/sync_rd[1]~FF .CE_POLARITY = 1'b1;
    defparam \fifo_inst/sync_rd[1]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/sync_rd[1]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/sync_rd[1]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/sync_rd[1]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/sync_rd[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[0][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[0][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[0][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[0][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[0][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[0][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[1][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[1][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[1][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[1][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[1][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[1][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[1][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[1][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[1][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[1][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[2][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[2][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[2][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[2][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[2][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[2][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[2][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[2][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[2][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[2][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[2][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[2][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[2][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[2][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[2][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[1]~FF  (.D(\fifo_inst/n143 ), .CE(ceg_net418), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/buff_head[1]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[1]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[1]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[1]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[1]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[1]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[2]~FF  (.D(\fifo_inst/n142 ), .CE(ceg_net418), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/buff_head[2]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[2]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[2]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[2]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[2]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[2]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[3]~FF  (.D(\fifo_inst/n141 ), .CE(ceg_net418), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/buff_head[3]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[3]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[3]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[3]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[3]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[3]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[4]~FF  (.D(\fifo_inst/n140 ), .CE(ceg_net418), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/buff_head[4]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[4]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[4]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[4]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[4]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[4]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[5]~FF  (.D(\fifo_inst/n139 ), .CE(ceg_net418), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/buff_head[5]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[5]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[5]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[5]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[5]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[5]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[6]~FF  (.D(\fifo_inst/n138 ), .CE(ceg_net418), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/buff_head[6]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[6]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[6]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[6]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[6]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[6]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \fifo_inst/buff_head[7]~FF  (.D(\fifo_inst/n137 ), .CE(ceg_net418), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\fifo_inst/buff_head[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \fifo_inst/buff_head[7]~FF .CLK_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[7]~FF .CE_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[7]~FF .SR_POLARITY = 1'b0;
    defparam \fifo_inst/buff_head[7]~FF .D_POLARITY = 1'b1;
    defparam \fifo_inst/buff_head[7]~FF .SR_SYNC = 1'b0;
    defparam \fifo_inst/buff_head[7]~FF .SR_VALUE = 1'b0;
    defparam \fifo_inst/buff_head[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/wr_index[0]~FF  (.D(\tx_fifo/n153 ), .CE(ceg_net234), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/wr_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/wr_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/wr_index[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/wr_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/rd_index[0]~FF  (.D(\tx_fifo/n162 ), .CE(ceg_net252), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/rd_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/rd_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/rd_index[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/rd_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/length[0]~FF  (.D(\data_to_tx_packet_len_reg[0] ), .CE(rx_en_tx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/length[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/length[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/length[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_fifo/length[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/length[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/length[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/length[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/length[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/sync_wr[0]~FF  (.D(rx_en_tx_packet), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\tx_fifo/sync_wr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/sync_wr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/sync_wr[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_fifo/sync_wr[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/sync_wr[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/sync_wr[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/sync_wr[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/sync_wr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/sync_rd[0]~FF  (.D(tx_en_tx_packet), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\tx_fifo/sync_rd[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/sync_rd[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/sync_rd[0]~FF .CE_POLARITY = 1'b1;
    defparam \tx_fifo/sync_rd[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/sync_rd[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/sync_rd[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/sync_rd[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/sync_rd[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/buff_head[0]~FF  (.D(\tx_fifo/n144 ), .CE(ceg_net458), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/buff_head[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/buff_head[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[0]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[0]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[0]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[0]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/buff_head[0]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/buff_head[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/wr_index[1]~FF  (.D(\tx_fifo/n152 ), .CE(ceg_net234), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/wr_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/wr_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/wr_index[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/wr_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/wr_index[2]~FF  (.D(\tx_fifo/n151 ), .CE(ceg_net234), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/wr_index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/wr_index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[2]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[2]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[2]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[2]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/wr_index[2]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/wr_index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/wr_index[3]~FF  (.D(\tx_fifo/n150 ), .CE(ceg_net234), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/wr_index[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/wr_index[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[3]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[3]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[3]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[3]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/wr_index[3]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/wr_index[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/wr_index[4]~FF  (.D(\tx_fifo/n149 ), .CE(ceg_net234), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/wr_index[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/wr_index[4]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[4]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[4]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[4]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[4]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/wr_index[4]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/wr_index[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/wr_index[5]~FF  (.D(\tx_fifo/n148 ), .CE(ceg_net234), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/wr_index[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/wr_index[5]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[5]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[5]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[5]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[5]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/wr_index[5]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/wr_index[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/wr_index[6]~FF  (.D(\tx_fifo/n147 ), .CE(ceg_net234), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/wr_index[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/wr_index[6]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[6]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[6]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[6]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[6]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/wr_index[6]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/wr_index[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/wr_index[7]~FF  (.D(\tx_fifo/n146 ), .CE(ceg_net234), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/wr_index[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/wr_index[7]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[7]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[7]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/wr_index[7]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/wr_index[7]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/wr_index[7]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/wr_index[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/rd_index[1]~FF  (.D(\tx_fifo/n161 ), .CE(ceg_net252), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/rd_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/rd_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/rd_index[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/rd_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/rd_index[2]~FF  (.D(\tx_fifo/n160 ), .CE(ceg_net252), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/rd_index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/rd_index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[2]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[2]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[2]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[2]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/rd_index[2]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/rd_index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/rd_index[3]~FF  (.D(\tx_fifo/n159 ), .CE(ceg_net252), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/rd_index[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/rd_index[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[3]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[3]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[3]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[3]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/rd_index[3]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/rd_index[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/rd_index[4]~FF  (.D(\tx_fifo/n158 ), .CE(ceg_net252), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/rd_index[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/rd_index[4]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[4]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[4]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[4]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[4]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/rd_index[4]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/rd_index[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/rd_index[5]~FF  (.D(\tx_fifo/n157 ), .CE(ceg_net252), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/rd_index[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/rd_index[5]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[5]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[5]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[5]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[5]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/rd_index[5]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/rd_index[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/rd_index[6]~FF  (.D(\tx_fifo/n156 ), .CE(ceg_net252), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/rd_index[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/rd_index[6]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[6]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[6]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[6]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[6]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/rd_index[6]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/rd_index[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/rd_index[7]~FF  (.D(\tx_fifo/n155 ), .CE(ceg_net252), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/rd_index[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/rd_index[7]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[7]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[7]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/rd_index[7]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/rd_index[7]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/rd_index[7]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/rd_index[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/length[1]~FF  (.D(\data_to_tx_packet_len_reg[1] ), .CE(rx_en_tx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/length[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/length[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/length[1]~FF .CE_POLARITY = 1'b1;
    defparam \tx_fifo/length[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/length[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/length[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/length[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/length[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/length[2]~FF  (.D(\data_to_tx_packet_len_reg[2] ), .CE(rx_en_tx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/length[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/length[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/length[2]~FF .CE_POLARITY = 1'b1;
    defparam \tx_fifo/length[2]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/length[2]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/length[2]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/length[2]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/length[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/length[3]~FF  (.D(\data_to_tx_packet_len_reg[3] ), .CE(rx_en_tx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/length[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/length[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/length[3]~FF .CE_POLARITY = 1'b1;
    defparam \tx_fifo/length[3]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/length[3]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/length[3]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/length[3]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/length[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/length[4]~FF  (.D(\data_to_tx_packet_len_reg[4] ), .CE(rx_en_tx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/length[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/length[4]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/length[4]~FF .CE_POLARITY = 1'b1;
    defparam \tx_fifo/length[4]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/length[4]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/length[4]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/length[4]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/length[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/length[5]~FF  (.D(\data_to_tx_packet_len_reg[5] ), .CE(rx_en_tx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/length[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/length[5]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/length[5]~FF .CE_POLARITY = 1'b1;
    defparam \tx_fifo/length[5]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/length[5]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/length[5]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/length[5]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/length[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/length[6]~FF  (.D(\data_to_tx_packet_len_reg[6] ), .CE(rx_en_tx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/length[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/length[6]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/length[6]~FF .CE_POLARITY = 1'b1;
    defparam \tx_fifo/length[6]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/length[6]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/length[6]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/length[6]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/length[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/length[7]~FF  (.D(\data_to_tx_packet_len_reg[7] ), .CE(rx_en_tx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/length[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/length[7]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/length[7]~FF .CE_POLARITY = 1'b1;
    defparam \tx_fifo/length[7]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/length[7]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/length[7]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/length[7]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/length[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/sync_wr[1]~FF  (.D(\tx_fifo/sync_wr[0] ), .CE(1'b1), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/sync_wr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/sync_wr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/sync_wr[1]~FF .CE_POLARITY = 1'b1;
    defparam \tx_fifo/sync_wr[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/sync_wr[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/sync_wr[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/sync_wr[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/sync_wr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/sync_rd[1]~FF  (.D(\tx_fifo/sync_rd[0] ), .CE(1'b1), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/sync_rd[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/sync_rd[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/sync_rd[1]~FF .CE_POLARITY = 1'b1;
    defparam \tx_fifo/sync_rd[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/sync_rd[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/sync_rd[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/sync_rd[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/sync_rd[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[0][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[0][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[0][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[0][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[0][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[0][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[1][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[1][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[1][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[1][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[1][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[1][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[1][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[1][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[1][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[1][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[1][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[1][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[1][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[1][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[1][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[2][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[2][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[2][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[2][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[2][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/buff_head[1]~FF  (.D(\tx_fifo/n143 ), .CE(ceg_net458), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/buff_head[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/buff_head[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[1]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[1]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[1]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[1]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/buff_head[1]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/buff_head[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/buff_head[2]~FF  (.D(\tx_fifo/n142 ), .CE(ceg_net458), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/buff_head[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/buff_head[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[2]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[2]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[2]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[2]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/buff_head[2]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/buff_head[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/buff_head[3]~FF  (.D(\tx_fifo/n141 ), .CE(ceg_net458), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/buff_head[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/buff_head[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[3]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[3]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[3]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[3]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/buff_head[3]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/buff_head[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/buff_head[4]~FF  (.D(\tx_fifo/n140 ), .CE(ceg_net458), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/buff_head[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/buff_head[4]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[4]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[4]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[4]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[4]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/buff_head[4]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/buff_head[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/buff_head[5]~FF  (.D(\tx_fifo/n139 ), .CE(ceg_net458), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/buff_head[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/buff_head[5]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[5]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[5]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[5]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[5]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/buff_head[5]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/buff_head[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/buff_head[6]~FF  (.D(\tx_fifo/n138 ), .CE(ceg_net458), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/buff_head[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/buff_head[6]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[6]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[6]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[6]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[6]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/buff_head[6]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/buff_head[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_fifo/buff_head[7]~FF  (.D(\tx_fifo/n137 ), .CE(ceg_net458), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\tx_fifo/buff_head[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \tx_fifo/buff_head[7]~FF .CLK_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[7]~FF .CE_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[7]~FF .SR_POLARITY = 1'b0;
    defparam \tx_fifo/buff_head[7]~FF .D_POLARITY = 1'b1;
    defparam \tx_fifo/buff_head[7]~FF .SR_SYNC = 1'b0;
    defparam \tx_fifo/buff_head[7]~FF .SR_VALUE = 1'b0;
    defparam \tx_fifo/buff_head[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/wr_index[0]~FF  (.D(\rx_fifo/n153 ), .CE(ceg_net322), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/wr_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/wr_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[0]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[0]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/wr_index[0]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/wr_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/rd_index[0]~FF  (.D(\rx_fifo/n162 ), .CE(ceg_net340), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/rd_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/rd_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[0]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[0]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/rd_index[0]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/rd_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/length[0]~FF  (.D(\data_to_rx_packet_len_reg[0] ), .CE(rx_en_rx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/length[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/length[0]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/length[0]~FF .CE_POLARITY = 1'b1;
    defparam \rx_fifo/length[0]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/length[0]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/length[0]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/length[0]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/length[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/sync_wr[0]~FF  (.D(rx_en_rx_packet), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_fifo/sync_wr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/sync_wr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/sync_wr[0]~FF .CE_POLARITY = 1'b1;
    defparam \rx_fifo/sync_wr[0]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/sync_wr[0]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/sync_wr[0]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/sync_wr[0]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/sync_wr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/sync_rd[0]~FF  (.D(n4269), .CE(1'b1), .CLK(\pll_clk~O ), 
           .SR(reset_n), .Q(\rx_fifo/sync_rd[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/sync_rd[0]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/sync_rd[0]~FF .CE_POLARITY = 1'b1;
    defparam \rx_fifo/sync_rd[0]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/sync_rd[0]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/sync_rd[0]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/sync_rd[0]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/sync_rd[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/buff_head[0]~FF  (.D(\rx_fifo/n144 ), .CE(ceg_net498), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/buff_head[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/buff_head[0]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[0]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[0]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[0]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[0]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/buff_head[0]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/buff_head[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/wr_index[1]~FF  (.D(\rx_fifo/n152 ), .CE(ceg_net322), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/wr_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/wr_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[1]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[1]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/wr_index[1]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/wr_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/wr_index[2]~FF  (.D(\rx_fifo/n151 ), .CE(ceg_net322), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/wr_index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/wr_index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[2]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[2]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[2]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[2]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/wr_index[2]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/wr_index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/wr_index[3]~FF  (.D(\rx_fifo/n150 ), .CE(ceg_net322), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/wr_index[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/wr_index[3]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[3]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[3]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[3]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[3]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/wr_index[3]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/wr_index[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/wr_index[4]~FF  (.D(\rx_fifo/n149 ), .CE(ceg_net322), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/wr_index[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/wr_index[4]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[4]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[4]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[4]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[4]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/wr_index[4]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/wr_index[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/wr_index[5]~FF  (.D(\rx_fifo/n148 ), .CE(ceg_net322), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/wr_index[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/wr_index[5]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[5]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[5]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[5]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[5]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/wr_index[5]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/wr_index[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/wr_index[6]~FF  (.D(\rx_fifo/n147 ), .CE(ceg_net322), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/wr_index[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/wr_index[6]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[6]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[6]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[6]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[6]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/wr_index[6]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/wr_index[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/wr_index[7]~FF  (.D(\rx_fifo/n146 ), .CE(ceg_net322), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/wr_index[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/wr_index[7]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[7]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[7]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/wr_index[7]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/wr_index[7]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/wr_index[7]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/wr_index[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/rd_index[1]~FF  (.D(\rx_fifo/n161 ), .CE(ceg_net340), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/rd_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/rd_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[1]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[1]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/rd_index[1]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/rd_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/rd_index[2]~FF  (.D(\rx_fifo/n160 ), .CE(ceg_net340), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/rd_index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/rd_index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[2]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[2]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[2]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[2]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/rd_index[2]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/rd_index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/rd_index[3]~FF  (.D(\rx_fifo/n159 ), .CE(ceg_net340), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/rd_index[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/rd_index[3]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[3]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[3]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[3]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[3]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/rd_index[3]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/rd_index[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/rd_index[4]~FF  (.D(\rx_fifo/n158 ), .CE(ceg_net340), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/rd_index[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/rd_index[4]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[4]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[4]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[4]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[4]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/rd_index[4]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/rd_index[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/rd_index[5]~FF  (.D(\rx_fifo/n157 ), .CE(ceg_net340), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/rd_index[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/rd_index[5]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[5]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[5]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[5]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[5]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/rd_index[5]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/rd_index[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/rd_index[6]~FF  (.D(\rx_fifo/n156 ), .CE(ceg_net340), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/rd_index[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/rd_index[6]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[6]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[6]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[6]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[6]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/rd_index[6]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/rd_index[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/rd_index[7]~FF  (.D(\rx_fifo/n155 ), .CE(ceg_net340), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/rd_index[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/rd_index[7]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[7]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[7]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/rd_index[7]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/rd_index[7]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/rd_index[7]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/rd_index[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/length[1]~FF  (.D(\data_to_rx_packet_len_reg[1] ), .CE(rx_en_rx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/length[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/length[1]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/length[1]~FF .CE_POLARITY = 1'b1;
    defparam \rx_fifo/length[1]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/length[1]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/length[1]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/length[1]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/length[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/length[2]~FF  (.D(\data_to_rx_packet_len_reg[2] ), .CE(rx_en_rx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/length[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/length[2]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/length[2]~FF .CE_POLARITY = 1'b1;
    defparam \rx_fifo/length[2]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/length[2]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/length[2]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/length[2]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/length[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/length[3]~FF  (.D(\data_to_rx_packet_len_reg[3] ), .CE(rx_en_rx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/length[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/length[3]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/length[3]~FF .CE_POLARITY = 1'b1;
    defparam \rx_fifo/length[3]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/length[3]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/length[3]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/length[3]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/length[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/length[4]~FF  (.D(\data_to_rx_packet_len_reg[4] ), .CE(rx_en_rx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/length[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/length[4]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/length[4]~FF .CE_POLARITY = 1'b1;
    defparam \rx_fifo/length[4]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/length[4]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/length[4]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/length[4]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/length[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/length[5]~FF  (.D(\data_to_rx_packet_len_reg[5] ), .CE(rx_en_rx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/length[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/length[5]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/length[5]~FF .CE_POLARITY = 1'b1;
    defparam \rx_fifo/length[5]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/length[5]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/length[5]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/length[5]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/length[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/length[6]~FF  (.D(\data_to_rx_packet_len_reg[6] ), .CE(rx_en_rx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/length[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/length[6]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/length[6]~FF .CE_POLARITY = 1'b1;
    defparam \rx_fifo/length[6]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/length[6]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/length[6]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/length[6]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/length[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/length[7]~FF  (.D(\data_to_rx_packet_len_reg[7] ), .CE(rx_en_rx_packet_len), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/length[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/length[7]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/length[7]~FF .CE_POLARITY = 1'b1;
    defparam \rx_fifo/length[7]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/length[7]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/length[7]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/length[7]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/length[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/sync_wr[1]~FF  (.D(\rx_fifo/sync_wr[0] ), .CE(1'b1), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/sync_wr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/sync_wr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/sync_wr[1]~FF .CE_POLARITY = 1'b1;
    defparam \rx_fifo/sync_wr[1]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/sync_wr[1]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/sync_wr[1]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/sync_wr[1]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/sync_wr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/sync_rd[1]~FF  (.D(\rx_fifo/sync_rd[0] ), .CE(1'b1), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/sync_rd[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/sync_rd[1]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/sync_rd[1]~FF .CE_POLARITY = 1'b1;
    defparam \rx_fifo/sync_rd[1]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/sync_rd[1]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/sync_rd[1]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/sync_rd[1]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/sync_rd[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[0][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[0][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[0][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[0][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[0][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[1][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[1][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[1][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[1][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[1][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[1][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[1][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[1][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[1][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[1][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[1][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[1][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[1][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[1][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[1][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[1][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[2][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[2][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[2][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[2][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[2][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[2][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[2][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[2][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[2][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[2][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[2][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/buff_head[1]~FF  (.D(\rx_fifo/n143 ), .CE(ceg_net498), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/buff_head[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/buff_head[1]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[1]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[1]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[1]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[1]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/buff_head[1]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/buff_head[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/buff_head[2]~FF  (.D(\rx_fifo/n142 ), .CE(ceg_net498), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/buff_head[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/buff_head[2]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[2]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[2]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[2]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[2]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/buff_head[2]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/buff_head[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/buff_head[3]~FF  (.D(\rx_fifo/n141 ), .CE(ceg_net498), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/buff_head[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/buff_head[3]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[3]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[3]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[3]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[3]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/buff_head[3]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/buff_head[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/buff_head[4]~FF  (.D(\rx_fifo/n140 ), .CE(ceg_net498), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/buff_head[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/buff_head[4]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[4]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[4]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[4]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[4]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/buff_head[4]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/buff_head[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/buff_head[5]~FF  (.D(\rx_fifo/n139 ), .CE(ceg_net498), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/buff_head[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/buff_head[5]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[5]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[5]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[5]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[5]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/buff_head[5]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/buff_head[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/buff_head[6]~FF  (.D(\rx_fifo/n138 ), .CE(ceg_net498), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/buff_head[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/buff_head[6]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[6]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[6]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[6]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[6]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/buff_head[6]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/buff_head[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rx_fifo/buff_head[7]~FF  (.D(\rx_fifo/n137 ), .CE(ceg_net498), 
           .CLK(\pll_clk~O ), .SR(reset_n), .Q(\rx_fifo/buff_head[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(76)
    defparam \rx_fifo/buff_head[7]~FF .CLK_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[7]~FF .CE_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[7]~FF .SR_POLARITY = 1'b0;
    defparam \rx_fifo/buff_head[7]~FF .D_POLARITY = 1'b1;
    defparam \rx_fifo/buff_head[7]~FF .SR_SYNC = 1'b0;
    defparam \rx_fifo/buff_head[7]~FF .SR_VALUE = 1'b0;
    defparam \rx_fifo/buff_head[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[3][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[3][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[3][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[3][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[3][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[3][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[3][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[3][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[3][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[3][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[3][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[3][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[3][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[3][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[3][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[3][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[3][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[3][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[3][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[3][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[3][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[3][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[3][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[3][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[3][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[3][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[4][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[4][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[4][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[4][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[4][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[4][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[4][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[4][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[4][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[4][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[4][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[4][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[4][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[4][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[4][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[4][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[4][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[4][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[4][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[4][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[4][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[4][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[4][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[4][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[4][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[4][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[4][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[4][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[4][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[4][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[4][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[4][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[4][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[4][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[4][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[4][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[4][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[4][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[4][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[4][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[4][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[5][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[5][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[5][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[5][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[5][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[5][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[5][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[5][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[5][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[5][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[5][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[5][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[5][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[5][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[5][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[5][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[5][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[5][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[5][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[5][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[5][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[5][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[5][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[5][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[5][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[5][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[5][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[5][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[5][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[5][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[5][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[5][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[5][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[5][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[5][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[5][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[5][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[5][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[5][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[5][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[5][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[6][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[6][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[6][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[6][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[6][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[6][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[6][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[6][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[6][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[6][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[6][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[6][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[6][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[6][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[6][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[6][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[6][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[6][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[6][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[6][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[6][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[6][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[6][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[6][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[6][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[6][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[6][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[6][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[6][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[6][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[6][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[6][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[6][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[6][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[6][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[6][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[6][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[6][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[6][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[6][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[6][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[7][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[7][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[7][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[7][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[7][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[7][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[7][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[7][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[7][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[7][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[7][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[7][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[7][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[7][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[7][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[7][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[7][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[7][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[7][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[7][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[7][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[7][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[7][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[7][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[7][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[7][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[7][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[7][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[7][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[7][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[7][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[7][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[7][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[7][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[7][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[7][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[7][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[7][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[7][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[7][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[7][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[8][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[8][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[8][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[8][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[8][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[8][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[8][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[8][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[8][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[8][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[8][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[8][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[8][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[8][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[8][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[8][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[8][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[8][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[8][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[8][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[8][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[8][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[8][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[8][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[8][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[8][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[8][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[8][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[8][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[8][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[8][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[8][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[8][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[8][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[8][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[8][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[8][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[8][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[8][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[8][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[8][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[9][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[9][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[9][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[9][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[9][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[9][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[9][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[9][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[9][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[9][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[9][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[9][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[9][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[9][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[9][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[9][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[9][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[9][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[9][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[9][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[9][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[9][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[9][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[9][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[9][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[9][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[9][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[9][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[9][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[9][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[9][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[9][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[9][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[9][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[9][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[9][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[9][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[9][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[9][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[9][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[9][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[10][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[10][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[10][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[10][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[10][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[10][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[10][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[10][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[10][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[10][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[10][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[10][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[10][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[10][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[10][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[10][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[10][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[10][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[10][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[10][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[10][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[10][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[10][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[10][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[10][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[10][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[10][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[10][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[10][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[10][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[10][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[10][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[10][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[10][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[10][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[10][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[10][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[10][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[10][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[10][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[10][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[11][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[11][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[11][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[11][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[11][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[11][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[11][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[11][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[11][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[11][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[11][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[11][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[11][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[11][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[11][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[11][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[11][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[11][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[11][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[11][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[11][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[11][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[11][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[11][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[11][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[11][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[11][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[11][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[11][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[11][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[11][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[11][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[11][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[11][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[11][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[11][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[11][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[11][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[11][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[11][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[11][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[12][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[12][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[12][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[12][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[12][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[12][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[12][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[12][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[12][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[12][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[12][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[12][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[12][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[12][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[12][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[12][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[12][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[12][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[12][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[12][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[12][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[12][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[12][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[12][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[12][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[12][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[12][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[12][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[12][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[12][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[12][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[12][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[12][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[12][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[12][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[12][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[12][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[12][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[12][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[12][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[12][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[13][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[13][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[13][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[13][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[13][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[13][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[13][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[13][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[13][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[13][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[13][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[13][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[13][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[13][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[13][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[13][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[13][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[13][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[13][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[13][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[13][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[13][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[13][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[13][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[13][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[13][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[13][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[13][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[13][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[13][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[13][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[13][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[13][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[13][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[13][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[13][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[13][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[13][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[13][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[13][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[13][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[14][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[14][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[14][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[14][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[14][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[14][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[14][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[14][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[14][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[14][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[14][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[14][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[14][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[14][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[14][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[14][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[14][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[14][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[14][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[14][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[14][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[14][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[14][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[14][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[14][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[14][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[14][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[14][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[14][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[14][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[14][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[14][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[14][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[14][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[14][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[14][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[14][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[14][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[14][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[14][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[14][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[15][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[15][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[15][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[15][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[15][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[15][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[15][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[15][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[15][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[15][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[15][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[15][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[15][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[15][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[15][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[15][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[15][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[15][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[15][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[15][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[15][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[15][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[15][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[15][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[15][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[15][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[15][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[15][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[15][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[15][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[15][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[15][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[15][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[15][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[15][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[15][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[15][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[15][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[15][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[15][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[15][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[16][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[16][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[16][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[16][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[16][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[16][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[16][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[16][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[16][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[16][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[16][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[16][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[16][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[16][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[16][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[16][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[16][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[16][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[16][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[16][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[16][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[16][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[16][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[16][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[16][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[16][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[16][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[16][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[16][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[16][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[16][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[16][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[16][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[16][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[16][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[16][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[16][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[16][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[16][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[16][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[16][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[17][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[17][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[17][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[17][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[17][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[17][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[17][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[17][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[17][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[17][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[17][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[17][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[17][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[17][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[17][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[17][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[17][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[17][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[17][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[17][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[17][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[17][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[17][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[17][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[17][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[17][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[17][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[17][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[17][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[17][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[17][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[17][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[17][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[17][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[17][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[17][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[17][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[17][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[17][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[17][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[17][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[18][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[18][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[18][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[18][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[18][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[18][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[18][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[18][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[18][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[18][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[18][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[18][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[18][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[18][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[18][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[18][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[18][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[18][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[18][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[18][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[18][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[18][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[18][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[18][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[18][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[18][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[18][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[18][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[18][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[18][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[18][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[18][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[18][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[18][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[18][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[18][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[18][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[18][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[18][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[18][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[18][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[19][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[19][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[19][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[19][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[19][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[19][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[19][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[19][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[19][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[19][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[19][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[19][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[19][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[19][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[19][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[19][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[19][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[19][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[19][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[19][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[19][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[19][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[19][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[19][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[19][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[19][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[19][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[19][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[19][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[19][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[19][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[19][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[19][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[19][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[19][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[19][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[19][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[19][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[19][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[19][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[19][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[20][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[20][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[20][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[20][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[20][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[20][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[20][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[20][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[20][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[20][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[20][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[20][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[20][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[20][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[20][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[20][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[20][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[20][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[20][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[20][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[20][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[20][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[20][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[20][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[20][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[20][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[20][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[20][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[20][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[20][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[20][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[20][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[20][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[20][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[20][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[20][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[20][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[20][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[20][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[20][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[20][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[21][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[21][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[21][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[21][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[21][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[21][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[21][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[21][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[21][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[21][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[21][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[21][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[21][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[21][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[21][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[21][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[21][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[21][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[21][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[21][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[21][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[21][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[21][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[21][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[21][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[21][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[21][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[21][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[21][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[21][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[21][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[21][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[21][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[21][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[21][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[21][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[21][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[21][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[21][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[21][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[21][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[22][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[22][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[22][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[22][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[22][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[22][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[22][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[22][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[22][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[22][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[22][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[22][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[22][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[22][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[22][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[22][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[22][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[22][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[22][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[22][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[22][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[22][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[22][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[22][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[22][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[22][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[22][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[22][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[22][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[22][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[22][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[22][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[22][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[22][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[22][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[22][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[22][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[22][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[22][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[22][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[22][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[23][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[23][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[23][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[23][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[23][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[23][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[23][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[23][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[23][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[23][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[23][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[23][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[23][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[23][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[23][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[23][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[23][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[23][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[23][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[23][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[23][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[23][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[23][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[23][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[23][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[23][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[23][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[23][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[23][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[23][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[23][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[23][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[23][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[23][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[23][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[23][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[23][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[23][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[23][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[23][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[23][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[24][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[24][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[24][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[24][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[24][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[24][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[24][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[24][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[24][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[24][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[24][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[24][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[24][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[24][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[24][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[24][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[24][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[24][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[24][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[24][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[24][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[24][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[24][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[24][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[24][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[24][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[24][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[24][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[24][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[24][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[24][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[24][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[24][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[24][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[24][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[24][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[24][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[24][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[24][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[24][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[24][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[25][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[25][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[25][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[25][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[25][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[25][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[25][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[25][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[25][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[25][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[25][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[25][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[25][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[25][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[25][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[25][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[25][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[25][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[25][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[25][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[25][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[25][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[25][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[25][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[25][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[25][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[25][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[25][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[25][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[25][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[25][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[25][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[25][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[25][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[25][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[25][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[25][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[25][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[25][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[25][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[25][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[26][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[26][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[26][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[26][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[26][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[26][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[26][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[26][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[26][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[26][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[26][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[26][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[26][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[26][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[26][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[26][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[26][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[26][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[26][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[26][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[26][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[26][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[26][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[26][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[26][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[26][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[26][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[26][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[26][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[26][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[26][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[26][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[26][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[26][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[26][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[26][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[26][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[26][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[26][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[26][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[26][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[27][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[27][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[27][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[27][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[27][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[27][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[27][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[27][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[27][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[27][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[27][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[27][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[27][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[27][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[27][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[27][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[27][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[27][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[27][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[27][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[27][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[27][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[27][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[27][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[27][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[27][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[27][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[27][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[27][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[27][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[27][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[27][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[27][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[27][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[27][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[27][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[27][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[27][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[27][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[27][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[27][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[28][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[28][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[28][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[28][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[28][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[28][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[28][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[28][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[28][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[28][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[28][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[28][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[28][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[28][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[28][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[28][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[28][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[28][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[28][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[28][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[28][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[28][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[28][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[28][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[28][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[28][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[28][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[28][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[28][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[28][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[28][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[28][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[28][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[28][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[28][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[28][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[28][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[28][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[28][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[28][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[28][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[29][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[29][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[29][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[29][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[29][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[29][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[29][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[29][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[29][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[29][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[29][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[29][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[29][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[29][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[29][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[29][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[29][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[29][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[29][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[29][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[29][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[29][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[29][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[29][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[29][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[29][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[29][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[29][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[29][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[29][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[29][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[29][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[29][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[29][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[29][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[29][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[29][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[29][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[29][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[29][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[29][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[30][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[30][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[30][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[30][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[30][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[30][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[30][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[30][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[30][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[30][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[30][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[30][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[30][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[30][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[30][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[30][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[30][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[30][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[30][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[30][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[30][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[30][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[30][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[30][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[30][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[30][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[30][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[30][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[30][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[30][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[30][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[30][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[30][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[30][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[30][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[30][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[30][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[30][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[30][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[30][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[30][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[31][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[31][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[31][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[31][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[31][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[31][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[31][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[31][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[31][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[31][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[31][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[31][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[31][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[31][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[31][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[31][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[31][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[31][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[31][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[31][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[31][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[31][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[31][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[31][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[31][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[31][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[31][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[31][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[31][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[31][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[31][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[31][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[31][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[31][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[31][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[31][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[31][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[31][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[31][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[31][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[31][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[32][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[32][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[32][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[32][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[32][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[32][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[32][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[32][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[32][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[32][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[32][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[32][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[32][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[32][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[32][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[32][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[32][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[32][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[32][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[32][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[32][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[32][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[32][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[32][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[32][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[32][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[32][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[32][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[32][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[32][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[32][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[32][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[32][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[32][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[32][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[32][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[32][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[32][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[32][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[32][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[32][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[33][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[33][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[33][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[33][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[33][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[33][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[33][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[33][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[33][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[33][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[33][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[33][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[33][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[33][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[33][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[33][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[33][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[33][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[33][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[33][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[33][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[33][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[33][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[33][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[33][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[33][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[33][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[33][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[33][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[33][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[33][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[33][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[33][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[33][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[33][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[33][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[33][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[33][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[33][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[33][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[33][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[34][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[34][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[34][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[34][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[34][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[34][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[34][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[34][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[34][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[34][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[34][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[34][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[34][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[34][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[34][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[34][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[34][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[34][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[34][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[34][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[34][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[34][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[34][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[34][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[34][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[34][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[34][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[34][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[34][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[34][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[34][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[34][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[34][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[34][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[34][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[34][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[34][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[34][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[34][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[34][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[34][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[35][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[35][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[35][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[35][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[35][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[35][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[35][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[35][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[35][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[35][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[35][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[35][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[35][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[35][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[35][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[35][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[35][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[35][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[35][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[35][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[35][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[35][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[35][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[35][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[35][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[35][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[35][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[35][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[35][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[35][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[35][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[35][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[35][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[35][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[35][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[35][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[35][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[35][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[35][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[35][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[35][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[36][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[36][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[36][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[36][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[36][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[36][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[36][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[36][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[36][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[36][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[36][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[36][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[36][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[36][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[36][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[36][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[36][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[36][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[36][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[36][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[36][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[36][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[36][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[36][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[36][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[36][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[36][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[36][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[36][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[36][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[36][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[36][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[36][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[36][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[36][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[36][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[36][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[36][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[36][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[36][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[36][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[37][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[37][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[37][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[37][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[37][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[37][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[37][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[37][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[37][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[37][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[37][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[37][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[37][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[37][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[37][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[37][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[37][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[37][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[37][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[37][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[37][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[37][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[37][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[37][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[37][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[37][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[37][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[37][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[37][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[37][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[37][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[37][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[37][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[37][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[37][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[37][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[37][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[37][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[37][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[37][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[37][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[38][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[38][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[38][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[38][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[38][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[38][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[38][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[38][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[38][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[38][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[38][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[38][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[38][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[38][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[38][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[38][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[38][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[38][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[38][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[38][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[38][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[38][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[38][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[38][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[38][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[38][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[38][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[38][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[38][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[38][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[38][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[38][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[38][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[38][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[38][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[38][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[38][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[38][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[38][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[38][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[38][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[39][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[39][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[39][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[39][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[39][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[39][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[39][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[39][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[39][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[39][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[39][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[39][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[39][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[39][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[39][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[39][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[39][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[39][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[39][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[39][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[39][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[39][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[39][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[39][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[39][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[39][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[39][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[39][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[39][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[39][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[39][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[39][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[39][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[39][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[39][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[39][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[39][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[39][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[39][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[39][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[39][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[40][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[40][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[40][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[40][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[40][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[40][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[40][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[40][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[40][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[40][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[40][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[40][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[40][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[40][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[40][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[40][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[40][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[40][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[40][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[40][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[40][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[40][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[40][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[40][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[40][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[40][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[40][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[40][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[40][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[40][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[40][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[40][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[40][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[40][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[40][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[40][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[40][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[40][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[40][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[40][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[40][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[41][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[41][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[41][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[41][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[41][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[41][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[41][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[41][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[41][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[41][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[41][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[41][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[41][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[41][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[41][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[41][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[41][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[41][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[41][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[41][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[41][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[41][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[41][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[41][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[41][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[41][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[41][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[41][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[41][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[41][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[41][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[41][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[41][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[41][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[41][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[41][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[41][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[41][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[41][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[41][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[41][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[42][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[42][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[42][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[42][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[42][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[42][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[42][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[42][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[42][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[42][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[42][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[42][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[42][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[42][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[42][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[42][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[42][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[42][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[42][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[42][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[42][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[42][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[42][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[42][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[42][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[42][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[42][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[42][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[42][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[42][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[42][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[42][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[42][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[42][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[42][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[42][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[42][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[42][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[42][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[42][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[42][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[43][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[43][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[43][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[43][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[43][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[43][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[43][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[43][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[43][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[43][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[43][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[43][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[43][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[43][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[43][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[43][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[43][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[43][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[43][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[43][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[43][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[43][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[43][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[43][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[43][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[43][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[43][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[43][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[43][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[43][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[43][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[43][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[43][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[43][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[43][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[43][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[43][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[43][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[43][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[43][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[43][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[44][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[44][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[44][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[44][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[44][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[44][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[44][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[44][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[44][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[44][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[44][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[44][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[44][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[44][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[44][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[44][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[44][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[44][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[44][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[44][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[44][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[44][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[44][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[44][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[44][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[44][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[44][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[44][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[44][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[44][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[44][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[44][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[44][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[44][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[44][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[44][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[44][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[44][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[44][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[44][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[44][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[45][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[45][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[45][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[45][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[45][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[45][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[45][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[45][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[45][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[45][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[45][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[45][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[45][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[45][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[45][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[45][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[45][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[45][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[45][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[45][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[45][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[45][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[45][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[45][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[45][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[45][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[45][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[45][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[45][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[45][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[45][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[45][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[45][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[45][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[45][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[45][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[45][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[45][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[45][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[45][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[45][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[46][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[46][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[46][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[46][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[46][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[46][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[46][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[46][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[46][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[46][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[46][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[46][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[46][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[46][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[46][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[46][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[46][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[46][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[46][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[46][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[46][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[46][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[46][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[46][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[46][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[46][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[46][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[46][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[46][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[46][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[46][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[46][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[46][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[46][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[46][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[46][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[46][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[46][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[46][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[46][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[46][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[47][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[47][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[47][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[47][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[47][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[47][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[47][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[47][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[47][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[47][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[47][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[47][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[47][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[47][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[47][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[47][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[47][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[47][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[47][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[47][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[47][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[47][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[47][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[47][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[47][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[47][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[47][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[47][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[47][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[47][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[47][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[47][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[47][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[47][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[47][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[47][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[47][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[47][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[47][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[47][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[47][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[48][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[48][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[48][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[48][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[48][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[48][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[48][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[48][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[48][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[48][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[48][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[48][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[48][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[48][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[48][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[48][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[48][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[48][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[48][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[48][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[48][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[48][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[48][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[48][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[48][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[48][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[48][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[48][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[48][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[48][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[48][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[48][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[48][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[48][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[48][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[48][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[48][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[48][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[48][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[48][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[48][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[49][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[49][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[49][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[49][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[49][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[49][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[49][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[49][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[49][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[49][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[49][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[49][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[49][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[49][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[49][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[49][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[49][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[49][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[49][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[49][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[49][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[49][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[49][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[49][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[49][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[49][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[49][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[49][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[49][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[49][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[49][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[49][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[49][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[49][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[49][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[49][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[49][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[49][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[49][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[49][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[49][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[50][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[50][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[50][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[50][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[50][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[50][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[50][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[50][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[50][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[50][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[50][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[50][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[50][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[50][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[50][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[50][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[50][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[50][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[50][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[50][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[50][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[50][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[50][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[50][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[50][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[50][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[50][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[50][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[50][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[50][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[50][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[50][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[50][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[50][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[50][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[50][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[50][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[50][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[50][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[50][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[50][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[51][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[51][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[51][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[51][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[51][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[51][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[51][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[51][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[51][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[51][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[51][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[51][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[51][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[51][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[51][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[51][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[51][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[51][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[51][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[51][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[51][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[51][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[51][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[51][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[51][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[51][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[51][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[51][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[51][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[51][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[51][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[51][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[51][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[51][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[51][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[51][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[51][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[51][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[51][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[51][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[51][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[52][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[52][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[52][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[52][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[52][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[52][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[52][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[52][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[52][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[52][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[52][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[52][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[52][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[52][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[52][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[52][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[52][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[52][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[52][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[52][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[52][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[52][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[52][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[52][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[52][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[52][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[52][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[52][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[52][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[52][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[52][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[52][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[52][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[52][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[52][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[52][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[52][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[52][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[52][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[52][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[52][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[53][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[53][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[53][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[53][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[53][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[53][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[53][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[53][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[53][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[53][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[53][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[53][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[53][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[53][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[53][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[53][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[53][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[53][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[53][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[53][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[53][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[53][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[53][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[53][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[53][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[53][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[53][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[53][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[53][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[53][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[53][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[53][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[53][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[53][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[53][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[53][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[53][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[53][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[53][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[53][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[53][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[54][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[54][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[54][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[54][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[54][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[54][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[54][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[54][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[54][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[54][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[54][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[54][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[54][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[54][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[54][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[54][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[54][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[54][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[54][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[54][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[54][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[54][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[54][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[54][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[54][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[54][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[54][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[54][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[54][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[54][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[54][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[54][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[54][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[54][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[54][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[54][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[54][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[54][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[54][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[54][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[54][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[55][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[55][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[55][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[55][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[55][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[55][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[55][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[55][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[55][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[55][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[55][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[55][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[55][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[55][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[55][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[55][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[55][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[55][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[55][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[55][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[55][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[55][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[55][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[55][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[55][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[55][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[55][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[55][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[55][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[55][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[55][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[55][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[55][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[55][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[55][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[55][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[55][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[55][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[55][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[55][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[55][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[56][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[56][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[56][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[56][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[56][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[56][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[56][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[56][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[56][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[56][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[56][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[56][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[56][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[56][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[56][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[56][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[56][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[56][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[56][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[56][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[56][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[56][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[56][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[56][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[56][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[56][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[56][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[56][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[56][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[56][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[56][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[56][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[56][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[56][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[56][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[56][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[56][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[56][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[56][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[56][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[56][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[57][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[57][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[57][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[57][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[57][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[57][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[57][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[57][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[57][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[57][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[57][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[57][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[57][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[57][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[57][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[57][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[57][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[57][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[57][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[57][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[57][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[57][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[57][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[57][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[57][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[57][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[57][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[57][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[57][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[57][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[57][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[57][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[57][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[57][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[57][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[57][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[57][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[57][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[57][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[57][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[57][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[58][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[58][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[58][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[58][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[58][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[58][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[58][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[58][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[58][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[58][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[58][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[58][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[58][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[58][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[58][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[58][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[58][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[58][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[58][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[58][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[58][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[58][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[58][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[58][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[58][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[58][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[58][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[58][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[58][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[58][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[58][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[58][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[58][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[58][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[58][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[58][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[58][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[58][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[58][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[58][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[58][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[59][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[59][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[59][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[59][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[59][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[59][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[59][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[59][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[59][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[59][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[59][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[59][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[59][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[59][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[59][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[59][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[59][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[59][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[59][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[59][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[59][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[59][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[59][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[59][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[59][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[59][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[59][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[59][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[59][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[59][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[59][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[59][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[59][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[59][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[59][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[59][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[59][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[59][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[59][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[59][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[59][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[60][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[60][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[60][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[60][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[60][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[60][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[60][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[60][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[60][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[60][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[60][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[60][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[60][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[60][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[60][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[60][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[60][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[60][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[60][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[60][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[60][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[60][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[60][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[60][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[60][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[60][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[60][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[60][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[60][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[60][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[60][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[60][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[60][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[60][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[60][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[60][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[60][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[60][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[60][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[60][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[60][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[61][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[61][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[61][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[61][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[61][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[61][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[61][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[61][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[61][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[61][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[61][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[61][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[61][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[61][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[61][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[61][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[61][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[61][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[61][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[61][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[61][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[61][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[61][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[61][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[61][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[61][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[61][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[61][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[61][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[61][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[61][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[61][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[61][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[61][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[61][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[61][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[61][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[61][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[61][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[61][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[61][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[62][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[62][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[62][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[62][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[62][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[62][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[62][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[62][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[62][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[62][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[62][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[62][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[62][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[62][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[62][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[62][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[62][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[62][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[62][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[62][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[62][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[62][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[62][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[62][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[62][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[62][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[62][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[62][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[62][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[62][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[62][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[62][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[62][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[62][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[62][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[62][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[62][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[62][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[62][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[62][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[62][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[63][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[63][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[63][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[63][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[63][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[63][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[63][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[63][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[63][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[63][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[63][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[63][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[63][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[63][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[63][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[63][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[63][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[63][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[63][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[63][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[63][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[63][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[63][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[63][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[63][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[63][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[63][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[63][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[63][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[63][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[63][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[63][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[63][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[63][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[63][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[63][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[63][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[63][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[63][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[63][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[63][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[64][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[64][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[64][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[64][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[64][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[64][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[64][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[64][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[64][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[64][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[64][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[64][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[64][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[64][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[64][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[64][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[64][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[64][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[64][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[64][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[64][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[64][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[64][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[64][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[64][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[64][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[64][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[64][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[64][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[64][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[64][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[64][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[64][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[64][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[64][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[64][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[64][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[64][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[64][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[64][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[64][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[65][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[65][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[65][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[65][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[65][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[65][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[65][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[65][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[65][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[65][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[65][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[65][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[65][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[65][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[65][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[65][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[65][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[65][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[65][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[65][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[65][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[65][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[65][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[65][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[65][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[65][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[65][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[65][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[65][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[65][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[65][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[65][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[65][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[65][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[65][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[65][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[65][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[65][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[65][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[65][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[65][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[66][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[66][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[66][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[66][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[66][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[66][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[66][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[66][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[66][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[66][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[66][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[66][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[66][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[66][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[66][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[66][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[66][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[66][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[66][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[66][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[66][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[66][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[66][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[66][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[66][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[66][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[66][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[66][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[66][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[66][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[66][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[66][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[66][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[66][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[66][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[66][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[66][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[66][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[66][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[66][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[66][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[67][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[67][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[67][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[67][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[67][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[67][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[67][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[67][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[67][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[67][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[67][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[67][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[67][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[67][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[67][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[67][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[67][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[67][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[67][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[67][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[67][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[67][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[67][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[67][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[67][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[67][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[67][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[67][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[67][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[67][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[67][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[67][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[67][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[67][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[67][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[67][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[67][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[67][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[67][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[67][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[67][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[68][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[68][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[68][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[68][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[68][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[68][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[68][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[68][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[68][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[68][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[68][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[68][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[68][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[68][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[68][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[68][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[68][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[68][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[68][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[68][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[68][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[68][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[68][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[68][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[68][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[68][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[68][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[68][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[68][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[68][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[68][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[68][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[68][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[68][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[68][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[68][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[68][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[68][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[68][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[68][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[68][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[69][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[69][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[69][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[69][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[69][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[69][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[69][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[69][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[69][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[69][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[69][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[69][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[69][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[69][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[69][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[69][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[69][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[69][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[69][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[69][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[69][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[69][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[69][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[69][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[69][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[69][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[69][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[69][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[69][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[69][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[69][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[69][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[69][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[69][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[69][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[69][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[69][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[69][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[69][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[69][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[69][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[70][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[70][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[70][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[70][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[70][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[70][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[70][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[70][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[70][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[70][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[70][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[70][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[70][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[70][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[70][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[70][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[70][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[70][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[70][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[70][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[70][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[70][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[70][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[70][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[70][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[70][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[70][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[70][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[70][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[70][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[70][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[70][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[70][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[70][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[70][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[70][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[70][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[70][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[70][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[70][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[70][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[71][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[71][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[71][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[71][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[71][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[71][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[71][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[71][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[71][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[71][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[71][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[71][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[71][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[71][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[71][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[71][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[71][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[71][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[71][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[71][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[71][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[71][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[71][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[71][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[71][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[71][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[71][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[71][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[71][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[71][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[71][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[71][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[71][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[71][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[71][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[71][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[71][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[71][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[71][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[71][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[71][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[72][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[72][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[72][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[72][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[72][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[72][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[72][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[72][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[72][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[72][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[72][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[72][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[72][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[72][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[72][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[72][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[72][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[72][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[72][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[72][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[72][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[72][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[72][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[72][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[72][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[72][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[72][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[72][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[72][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[72][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[72][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[72][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[72][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[72][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[72][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[72][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[72][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[72][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[72][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[72][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[72][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[73][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[73][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[73][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[73][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[73][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[73][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[73][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[73][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[73][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[73][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[73][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[73][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[73][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[73][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[73][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[73][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[73][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[73][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[73][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[73][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[73][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[73][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[73][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[73][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[73][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[73][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[73][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[73][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[73][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[73][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[73][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[73][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[73][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[73][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[73][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[73][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[73][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[73][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[73][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[73][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[73][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[74][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[74][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[74][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[74][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[74][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[74][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[74][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[74][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[74][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[74][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[74][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[74][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[74][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[74][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[74][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[74][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[74][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[74][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[74][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[74][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[74][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[74][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[74][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[74][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[74][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[74][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[74][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[74][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[74][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[74][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[74][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[74][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[74][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[74][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[74][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[74][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[74][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[74][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[74][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[74][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[74][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[75][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[75][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[75][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[75][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[75][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[75][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[75][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[75][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[75][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[75][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[75][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[75][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[75][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[75][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[75][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[75][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[75][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[75][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[75][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[75][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[75][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[75][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[75][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[75][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[75][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[75][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[75][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[75][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[75][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[75][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[75][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[75][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[75][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[75][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[75][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[75][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[75][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[75][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[75][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[75][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[75][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[76][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[76][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[76][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[76][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[76][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[76][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[76][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[76][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[76][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[76][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[76][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[76][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[76][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[76][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[76][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[76][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[76][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[76][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[76][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[76][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[76][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[76][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[76][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[76][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[76][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[76][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[76][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[76][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[76][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[76][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[76][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[76][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[76][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[76][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[76][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[76][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[76][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[76][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[76][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[76][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[76][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[77][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[77][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[77][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[77][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[77][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[77][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[77][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[77][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[77][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[77][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[77][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[77][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[77][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[77][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[77][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[77][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[77][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[77][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[77][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[77][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[77][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[77][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[77][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[77][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[77][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[77][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[77][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[77][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[77][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[77][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[77][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[77][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[77][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[77][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[77][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[77][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[77][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[77][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[77][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[77][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[77][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[78][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[78][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[78][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[78][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[78][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[78][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[78][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[78][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[78][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[78][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[78][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[78][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[78][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[78][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[78][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[78][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[78][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[78][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[78][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[78][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[78][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[78][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[78][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[78][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[78][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[78][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[78][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[78][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[78][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[78][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[78][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[78][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[78][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[78][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[78][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[78][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[78][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[78][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[78][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[78][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[78][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[79][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[79][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[79][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[79][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[79][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[79][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[79][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[79][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[79][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[79][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[79][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[79][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[79][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[79][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[79][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[79][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[79][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[79][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[79][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[79][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[79][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[79][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[79][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[79][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[79][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[79][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[79][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[79][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[79][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[79][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[79][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[79][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[79][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[79][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[79][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[79][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[79][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[79][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[79][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[79][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[79][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[80][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[80][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[80][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[80][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[80][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[80][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[80][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[80][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[80][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[80][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[80][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[80][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[80][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[80][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[80][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[80][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[80][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[80][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[80][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[80][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[80][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[80][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[80][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[80][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[80][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[80][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[80][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[80][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[80][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[80][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[80][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[80][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[80][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[80][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[80][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[80][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[80][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[80][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[80][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[80][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[80][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[81][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[81][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[81][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[81][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[81][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[81][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[81][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[81][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[81][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[81][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[81][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[81][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[81][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[81][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[81][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[81][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[81][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[81][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[81][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[81][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[81][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[81][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[81][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[81][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[81][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[81][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[81][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[81][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[81][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[81][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[81][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[81][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[81][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[81][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[81][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[81][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[81][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[81][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[81][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[81][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[81][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[82][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[82][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[82][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[82][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[82][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[82][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[82][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[82][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[82][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[82][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[82][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[82][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[82][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[82][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[82][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[82][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[82][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[82][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[82][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[82][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[82][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[82][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[82][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[82][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[82][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[82][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[82][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[82][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[82][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[82][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[82][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[82][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[82][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[82][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[82][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[82][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[82][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[82][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[82][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[82][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[82][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[83][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[83][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[83][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[83][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[83][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[83][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[83][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[83][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[83][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[83][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[83][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[83][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[83][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[83][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[83][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[83][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[83][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[83][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[83][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[83][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[83][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[83][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[83][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[83][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[83][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[83][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[83][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[83][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[83][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[83][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[83][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[83][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[83][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[83][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[83][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[83][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[83][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[83][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[83][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[83][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[83][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[84][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[84][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[84][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[84][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[84][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[84][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[84][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[84][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[84][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[84][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[84][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[84][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[84][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[84][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[84][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[84][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[84][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[84][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[84][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[84][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[84][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[84][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[84][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[84][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[84][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[84][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[84][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[84][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[84][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[84][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[84][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[84][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[84][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[84][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[84][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[84][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[84][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[84][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[84][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[84][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[84][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[85][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[85][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[85][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[85][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[85][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[85][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[85][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[85][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[85][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[85][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[85][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[85][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[85][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[85][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[85][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[85][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[85][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[85][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[85][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[85][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[85][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[85][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[85][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[85][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[85][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[85][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[85][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[85][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[85][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[85][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[85][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[85][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[85][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[85][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[85][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[85][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[85][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[85][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[85][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[85][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[85][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[86][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[86][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[86][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[86][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[86][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[86][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[86][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[86][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[86][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[86][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[86][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[86][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[86][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[86][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[86][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[86][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[86][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[86][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[86][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[86][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[86][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[86][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[86][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[86][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[86][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[86][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[86][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[86][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[86][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[86][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[86][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[86][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[86][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[86][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[86][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[86][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[86][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[86][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[86][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[86][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[86][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[87][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[87][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[87][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[87][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[87][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[87][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[87][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[87][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[87][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[87][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[87][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[87][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[87][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[87][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[87][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[87][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[87][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[87][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[87][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[87][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[87][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[87][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[87][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[87][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[87][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[87][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[87][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[87][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[87][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[87][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[87][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[87][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[87][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[87][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[87][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[87][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[87][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[87][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[87][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[87][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[87][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[88][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[88][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[88][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[88][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[88][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[88][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[88][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[88][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[88][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[88][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[88][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[88][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[88][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[88][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[88][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[88][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[88][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[88][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[88][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[88][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[88][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[88][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[88][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[88][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[88][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[88][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[88][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[88][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[88][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[88][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[88][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[88][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[88][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[88][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[88][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[88][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[88][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[88][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[88][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[88][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[88][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[89][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[89][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[89][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[89][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[89][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[89][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[89][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[89][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[89][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[89][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[89][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[89][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[89][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[89][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[89][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[89][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[89][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[89][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[89][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[89][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[89][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[89][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[89][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[89][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[89][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[89][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[89][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[89][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[89][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[89][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[89][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[89][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[89][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[89][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[89][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[89][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[89][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[89][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[89][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[89][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[89][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[90][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[90][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[90][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[90][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[90][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[90][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[90][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[90][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[90][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[90][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[90][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[90][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[90][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[90][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[90][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[90][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[90][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[90][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[90][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[90][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[90][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[90][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[90][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[90][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[90][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[90][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[90][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[90][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[90][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[90][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[90][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[90][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[90][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[90][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[90][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[90][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[90][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[90][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[90][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[90][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[90][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[91][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[91][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[91][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[91][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[91][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[91][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[91][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[91][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[91][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[91][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[91][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[91][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[91][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[91][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[91][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[91][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[91][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[91][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[91][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[91][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[91][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[91][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[91][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[91][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[91][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[91][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[91][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[91][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[91][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[91][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[91][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[91][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[91][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[91][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[91][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[91][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[91][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[91][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[91][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[91][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[91][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[92][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[92][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[92][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[92][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[92][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[92][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[92][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[92][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[92][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[92][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[92][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[92][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[92][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[92][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[92][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[92][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[92][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[92][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[92][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[92][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[92][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[92][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[92][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[92][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[92][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[92][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[92][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[92][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[92][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[92][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[92][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[92][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[92][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[92][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[92][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[92][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[92][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[92][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[92][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[92][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[92][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[93][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[93][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[93][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[93][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[93][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[93][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[93][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[93][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[93][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[93][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[93][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[93][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[93][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[93][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[93][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[93][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[93][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[93][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[93][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[93][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[93][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[93][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[93][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[93][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[93][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[93][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[93][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[93][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[93][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[93][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[93][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[93][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[93][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[93][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[93][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[93][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[93][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[93][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[93][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[93][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[93][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[94][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[94][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[94][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[94][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[94][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[94][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[94][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[94][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[94][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[94][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[94][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[94][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[94][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[94][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[94][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[94][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[94][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[94][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[94][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[94][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[94][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[94][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[94][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[94][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[94][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[94][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[94][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[94][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[94][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[94][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[94][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[94][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[94][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[94][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[94][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[94][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[94][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[94][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[94][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[94][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[94][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[95][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[95][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[95][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[95][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[95][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[95][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[95][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[95][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[95][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[95][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[95][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[95][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[95][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[95][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[95][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[95][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[95][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[95][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[95][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[95][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[95][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[95][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[95][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[95][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[95][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[95][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[95][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[95][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[95][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[95][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[95][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[95][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[95][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[95][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[95][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[95][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[95][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[95][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[95][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[95][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[95][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[96][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[96][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[96][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[96][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[96][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[96][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[96][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[96][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[96][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[96][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[96][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[96][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[96][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[96][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[96][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[96][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[96][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[96][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[96][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[96][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[96][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[96][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[96][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[96][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[96][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[96][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[96][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[96][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[96][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[96][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[96][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[96][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[96][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[96][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[96][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[96][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[96][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[96][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[96][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[96][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[96][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[97][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[97][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[97][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[97][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[97][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[97][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[97][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[97][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[97][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[97][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[97][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[97][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[97][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[97][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[97][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[97][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[97][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[97][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[97][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[97][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[97][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[97][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[97][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[97][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[97][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[97][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[97][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[97][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[97][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[97][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[97][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[97][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[97][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[97][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[97][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[97][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[97][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[97][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[97][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[97][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[97][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[98][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[98][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[98][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[98][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[98][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[98][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[98][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[98][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[98][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[98][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[98][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[98][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[98][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[98][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[98][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[98][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[98][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[98][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[98][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[98][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[98][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[98][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[98][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[98][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[98][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[98][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[98][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[98][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[98][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[98][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[98][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[98][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[98][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[98][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[98][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[98][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[98][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[98][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[98][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[98][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[98][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[99][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[99][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[99][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[99][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[99][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[99][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[99][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[99][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[99][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[99][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[99][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[99][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[99][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[99][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[99][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[99][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[99][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[99][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[99][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[99][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[99][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[99][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[99][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[99][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[99][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[99][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[99][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[99][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[99][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[99][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[99][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[99][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[99][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[99][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[99][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[99][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[99][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[99][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[99][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[99][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[99][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[100][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[100][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[100][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[100][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[100][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[100][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[100][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[100][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[100][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[100][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[100][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[100][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[100][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[100][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[100][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[100][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[100][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[100][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[100][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[100][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[100][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[100][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[100][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[100][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[100][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[100][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[100][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[100][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[100][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[100][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[100][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[100][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[100][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[100][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[100][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[100][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n32 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[100][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[100][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[100][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[100][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[100][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[101][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[101][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[101][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[101][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[101][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[101][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[101][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[101][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[101][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[101][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[101][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[101][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[101][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[101][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[101][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[101][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[101][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[101][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[101][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[101][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[101][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[101][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[101][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[101][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[101][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[101][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[101][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[101][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[101][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[101][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[101][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[101][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[101][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[101][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[101][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[101][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n31 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[101][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[101][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[101][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[101][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[101][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[102][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[102][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[102][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[102][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[102][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[102][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[102][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[102][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[102][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[102][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[102][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[102][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[102][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[102][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[102][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[102][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[102][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[102][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[102][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[102][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[102][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[102][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[102][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[102][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[102][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[102][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[102][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[102][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[102][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[102][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[102][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[102][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[102][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[102][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[102][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[102][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n30 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[102][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[102][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[102][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[102][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[102][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[103][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[103][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[103][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[103][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[103][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[103][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[103][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[103][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[103][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[103][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[103][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[103][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[103][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[103][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[103][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[103][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[103][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[103][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[103][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[103][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[103][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[103][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[103][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[103][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[103][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[103][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[103][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[103][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[103][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[103][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[103][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[103][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[103][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[103][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[103][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[103][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n29 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[103][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[103][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[103][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[103][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[103][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[104][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[104][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[104][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[104][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[104][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[104][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[104][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[104][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[104][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[104][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[104][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[104][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[104][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[104][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[104][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[104][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[104][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[104][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[104][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[104][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[104][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[104][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[104][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[104][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[104][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[104][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[104][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[104][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[104][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[104][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[104][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[104][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[104][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[104][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[104][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[104][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n28 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[104][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[104][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[104][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[104][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[104][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[105][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[105][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[105][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[105][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[105][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[105][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[105][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[105][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[105][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[105][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[105][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[105][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[105][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[105][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[105][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[105][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[105][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[105][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[105][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[105][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[105][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[105][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[105][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[105][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[105][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[105][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[105][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[105][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[105][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[105][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[105][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[105][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[105][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[105][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[105][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[105][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n27 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[105][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[105][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[105][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[105][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[105][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[106][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[106][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[106][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[106][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[106][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[106][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[106][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[106][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[106][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[106][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[106][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[106][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[106][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[106][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[106][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[106][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[106][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[106][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[106][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[106][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[106][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[106][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[106][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[106][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[106][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[106][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[106][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[106][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[106][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[106][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[106][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[106][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[106][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[106][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[106][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[106][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n26 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[106][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[106][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[106][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[106][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[106][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[107][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[107][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[107][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[107][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[107][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[107][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[107][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[107][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[107][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[107][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[107][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[107][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[107][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[107][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[107][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[107][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[107][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[107][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[107][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[107][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[107][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[107][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[107][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[107][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[107][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[107][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[107][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[107][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[107][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[107][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[107][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[107][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[107][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[107][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[107][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[107][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n25 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[107][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[107][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[107][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[107][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[107][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[108][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[108][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[108][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[108][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[108][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[108][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[108][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[108][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[108][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[108][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[108][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[108][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[108][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[108][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[108][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[108][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[108][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[108][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[108][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[108][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[108][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[108][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[108][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[108][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[108][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[108][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[108][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[108][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[108][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[108][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[108][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[108][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[108][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[108][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[108][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[108][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n24 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[108][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[108][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[108][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[108][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[108][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[109][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[109][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[109][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[109][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[109][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[109][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[109][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[109][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[109][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[109][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[109][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[109][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[109][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[109][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[109][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[109][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[109][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[109][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[109][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[109][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[109][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[109][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[109][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[109][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[109][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[109][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[109][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[109][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[109][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[109][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[109][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[109][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[109][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[109][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[109][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[109][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n23 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[109][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[109][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[109][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[109][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[109][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[110][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[110][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[110][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[110][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[110][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[110][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[110][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[110][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[110][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[110][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[110][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[110][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[110][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[110][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[110][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[110][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[110][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[110][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[110][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[110][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[110][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[110][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[110][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[110][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[110][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[110][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[110][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[110][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[110][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[110][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[110][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[110][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[110][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[110][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[110][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[110][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n22 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[110][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[110][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[110][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[110][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[110][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[111][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[111][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[111][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[111][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[111][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[111][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[111][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[111][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[111][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[111][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[111][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[111][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[111][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[111][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[111][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[111][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[111][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[111][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[111][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[111][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[111][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[111][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[111][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[111][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[111][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[111][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[111][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[111][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[111][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[111][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[111][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[111][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[111][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[111][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[111][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[111][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n21 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[111][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[111][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[111][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[111][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[111][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[112][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[112][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[112][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[112][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[112][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[112][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[112][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[112][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[112][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[112][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[112][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[112][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[112][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[112][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[112][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[112][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[112][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[112][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[112][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[112][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[112][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[112][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[112][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[112][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[112][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[112][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[112][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[112][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[112][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[112][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[112][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[112][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[112][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[112][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[112][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[112][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n20 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[112][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[112][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[112][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[112][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[112][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[113][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[113][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[113][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[113][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[113][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[113][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[113][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[113][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[113][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[113][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[113][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[113][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[113][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[113][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[113][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[113][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[113][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[113][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[113][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[113][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[113][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[113][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[113][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[113][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[113][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[113][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[113][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[113][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[113][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[113][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[113][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[113][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[113][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[113][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[113][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[113][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n19 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[113][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[113][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[113][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[113][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[113][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[114][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[114][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[114][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[114][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[114][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[114][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[114][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[114][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[114][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[114][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[114][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[114][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[114][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[114][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[114][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[114][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[114][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[114][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[114][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[114][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[114][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[114][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[114][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[114][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[114][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[114][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[114][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[114][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[114][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[114][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[114][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[114][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[114][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[114][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[114][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[114][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n18 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[114][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[114][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[114][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[114][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[114][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[115][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[115][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[115][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[115][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[115][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[115][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[115][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[115][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[115][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[115][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[115][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[115][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[115][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[115][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[115][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[115][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[115][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[115][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[115][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[115][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[115][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[115][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[115][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[115][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[115][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[115][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[115][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[115][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[115][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[115][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[115][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[115][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[115][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[115][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[115][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[115][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n17 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[115][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[115][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[115][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[115][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[115][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[116][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[116][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[116][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[116][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[116][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[116][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[116][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[116][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[116][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[116][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[116][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[116][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[116][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[116][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[116][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[116][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[116][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[116][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[116][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[116][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[116][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[116][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[116][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[116][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[116][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[116][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[116][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[116][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[116][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[116][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[116][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[116][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[116][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[116][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[116][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[116][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n16 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[116][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[116][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[116][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[116][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[116][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[117][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[117][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[117][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[117][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[117][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[117][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[117][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[117][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[117][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[117][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[117][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[117][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[117][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[117][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[117][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[117][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[117][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[117][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[117][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[117][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[117][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[117][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[117][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[117][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[117][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[117][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[117][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[117][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[117][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[117][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[117][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[117][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[117][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[117][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[117][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[117][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n15 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[117][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[117][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[117][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[117][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[117][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[118][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[118][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[118][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[118][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[118][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[118][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[118][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[118][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[118][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[118][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[118][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[118][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[118][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[118][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[118][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[118][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[118][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[118][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[118][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[118][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[118][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[118][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[118][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[118][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[118][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[118][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[118][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[118][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[118][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[118][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[118][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[118][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[118][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[118][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[118][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[118][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n14 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[118][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[118][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[118][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[118][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[118][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[119][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[119][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[119][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[119][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[119][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[119][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[119][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[119][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[119][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[119][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[119][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[119][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[119][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[119][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[119][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[119][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[119][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[119][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[119][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[119][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[119][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[119][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[119][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[119][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[119][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[119][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[119][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[119][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[119][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[119][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[119][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[119][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[119][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[119][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[119][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[119][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n13 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[119][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[119][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[119][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[119][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[119][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[120][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[120][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[120][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[120][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[120][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[120][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[120][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[120][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[120][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[120][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[120][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[120][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[120][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[120][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[120][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[120][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[120][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[120][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[120][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[120][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[120][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[120][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[120][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[120][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[120][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[120][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[120][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[120][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[120][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[120][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[120][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[120][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[120][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[120][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[120][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[120][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n12 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[120][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[120][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[120][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[120][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[120][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[121][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[121][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[121][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[121][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[121][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[121][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[121][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[121][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[121][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[121][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[121][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[121][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[121][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[121][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[121][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[121][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[121][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[121][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[121][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[121][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[121][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[121][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[121][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[121][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[121][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[121][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[121][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[121][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[121][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[121][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[121][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[121][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[121][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[121][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[121][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[121][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n11 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[121][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[121][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[121][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[121][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[121][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[122][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[122][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[122][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[122][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[122][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[122][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[122][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[122][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[122][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[122][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[122][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[122][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[122][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[122][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[122][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[122][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[122][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[122][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[122][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[122][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[122][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[122][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[122][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[122][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[122][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[122][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[122][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[122][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[122][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[122][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[122][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[122][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[122][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[122][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[122][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[122][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n10 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[122][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[122][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[122][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[122][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[122][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[123][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[123][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[123][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[123][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[123][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[123][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[123][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[123][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[123][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[123][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[123][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[123][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[123][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[123][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[123][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[123][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[123][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[123][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[123][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[123][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[123][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[123][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[123][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[123][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[123][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[123][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[123][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[123][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[123][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[123][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[123][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[123][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[123][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[123][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[123][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[123][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n9 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[123][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[123][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[123][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[123][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[123][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[124][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[124][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[124][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[124][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[124][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[124][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[124][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[124][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[124][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[124][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[124][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[124][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[124][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[124][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[124][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[124][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[124][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[124][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[124][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[124][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[124][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[124][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[124][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[124][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[124][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[124][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[124][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[124][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[124][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[124][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[124][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[124][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[124][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[124][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[124][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[124][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n8 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[124][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[124][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[124][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[124][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[124][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[125][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[125][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[125][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[125][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[125][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[125][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[125][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[125][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[125][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[125][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[125][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[125][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[125][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[125][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[125][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[125][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[125][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[125][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[125][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[125][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[125][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[125][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[125][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[125][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[125][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[125][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[125][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[125][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[125][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[125][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[125][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[125][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[125][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[125][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[125][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[125][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n7 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[125][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[125][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[125][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[125][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[125][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[126][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[126][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[126][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[126][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[126][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[126][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[126][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[126][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[126][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[126][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[126][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[126][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[126][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[126][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[126][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[126][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[126][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[126][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[126][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[126][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[126][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[126][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[126][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[126][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[126][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[126][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[126][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[126][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[126][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[126][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[126][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[126][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[126][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[126][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[126][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[126][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n6 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[126][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[126][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[126][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[126][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[126][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[127][0]~FF  (.D(\data_to_fifo[0] ), .CE(\i14/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[127][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[127][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][0]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][0]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][0]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][0]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[127][0]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[127][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[127][1]~FF  (.D(\data_to_fifo[1] ), .CE(\i14/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[127][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[127][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][1]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][1]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][1]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][1]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[127][1]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[127][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[127][2]~FF  (.D(\data_to_fifo[2] ), .CE(\i14/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[127][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[127][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][2]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][2]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][2]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][2]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[127][2]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[127][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[127][3]~FF  (.D(\data_to_fifo[3] ), .CE(\i14/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[127][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[127][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][3]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][3]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][3]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][3]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[127][3]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[127][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[127][4]~FF  (.D(\data_to_fifo[4] ), .CE(\i14/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[127][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[127][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][4]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][4]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][4]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][4]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[127][4]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[127][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[127][5]~FF  (.D(\data_to_fifo[5] ), .CE(\i14/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[127][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[127][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][5]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][5]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][5]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][5]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[127][5]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[127][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[127][6]~FF  (.D(\data_to_fifo[6] ), .CE(\i14/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[127][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[127][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][6]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][6]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][6]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][6]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[127][6]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[127][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i14/fifo_inst/buff[127][7]~FF  (.D(\data_to_fifo[7] ), .CE(\i14/n5 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i14/fifo_inst/buff[127][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i14/fifo_inst/buff[127][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][7]~FF .CE_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][7]~FF .SR_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][7]~FF .D_POLARITY = 1'b1;
    defparam \i14/fifo_inst/buff[127][7]~FF .SR_SYNC = 1'b1;
    defparam \i14/fifo_inst/buff[127][7]~FF .SR_VALUE = 1'b0;
    defparam \i14/fifo_inst/buff[127][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[0][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[0][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[0][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[0][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[0][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[0][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[0][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[0][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[0][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[0][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[0][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[0][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[0][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[0][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[0][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[0][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[0][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[1][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[1][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[1][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[1][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[1][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[1][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[1][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[1][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[1][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[1][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[1][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[1][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[1][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[1][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[1][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[1][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[1][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[1][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[1][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[1][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[1][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[1][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[1][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[1][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[1][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[1][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[1][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[1][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[1][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[1][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[1][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[1][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[1][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[1][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[1][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[1][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[1][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[1][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[1][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[1][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[1][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[2][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[2][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[2][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[2][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[2][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[2][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[2][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[2][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[2][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[2][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[2][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[2][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[2][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[2][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[2][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[2][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[2][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[2][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[2][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[2][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[2][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[2][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[2][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[2][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[2][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[2][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[2][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[2][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[2][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[2][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[2][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[2][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[2][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[2][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[2][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[2][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[2][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[2][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[2][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[2][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[2][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[3][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[3][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[3][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[3][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[3][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[3][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[3][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[3][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[3][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[3][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[3][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[3][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[3][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[3][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[3][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[3][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[3][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[3][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[3][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[3][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[3][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[3][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[3][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[3][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[3][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[3][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[3][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[3][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[3][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[3][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[3][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[3][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[3][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[3][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[3][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[3][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[3][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[3][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[3][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[3][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[3][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[4][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[4][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[4][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[4][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[4][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[4][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[4][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[4][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[4][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[4][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[4][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[4][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[4][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[4][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[4][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[4][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[4][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[4][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[4][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[4][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[4][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[4][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[4][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[4][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[4][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[4][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[4][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[4][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[4][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[4][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[4][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[4][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[4][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[4][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[4][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[4][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[4][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[4][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[4][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[4][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[4][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[5][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[5][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[5][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[5][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[5][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[5][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[5][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[5][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[5][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[5][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[5][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[5][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[5][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[5][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[5][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[5][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[5][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[5][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[5][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[5][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[5][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[5][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[5][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[5][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[5][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[5][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[5][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[5][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[5][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[5][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[5][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[5][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[5][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[5][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[5][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[5][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[5][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[5][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[5][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[5][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[5][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[6][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[6][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[6][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[6][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[6][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[6][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[6][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[6][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[6][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[6][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[6][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[6][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[6][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[6][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[6][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[6][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[6][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[6][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[6][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[6][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[6][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[6][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[6][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[6][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[6][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[6][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[6][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[6][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[6][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[6][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[6][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[6][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[6][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[6][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[6][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[6][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[6][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[6][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[6][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[6][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[6][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[7][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[7][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[7][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[7][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[7][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[7][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[7][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[7][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[7][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[7][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[7][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[7][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[7][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[7][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[7][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[7][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[7][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[7][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[7][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[7][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[7][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[7][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[7][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[7][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[7][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[7][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[7][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[7][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[7][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[7][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[7][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[7][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[7][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[7][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[7][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[7][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[7][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[7][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[7][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[7][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[7][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[8][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[8][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[8][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[8][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[8][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[8][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[8][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[8][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[8][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[8][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[8][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[8][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[8][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[8][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[8][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[8][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[8][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[8][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[8][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[8][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[8][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[8][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[8][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[8][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[8][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[8][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[8][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[8][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[8][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[8][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[8][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[8][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[8][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[8][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[8][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[8][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[8][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[8][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[8][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[8][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[8][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[9][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[9][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[9][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[9][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[9][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[9][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[9][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[9][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[9][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[9][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[9][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[9][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[9][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[9][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[9][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[9][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[9][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[9][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[9][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[9][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[9][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[9][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[9][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[9][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[9][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[9][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[9][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[9][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[9][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[9][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[9][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[9][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[9][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[9][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[9][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[9][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[9][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[9][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[9][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[9][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[9][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[10][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[10][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[10][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[10][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[10][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[10][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[10][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[10][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[10][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[10][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[10][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[10][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[10][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[10][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[10][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[10][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[10][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[10][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[10][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[10][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[10][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[10][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[10][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[10][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[10][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[10][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[10][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[10][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[10][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[10][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[10][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[10][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[10][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[10][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[10][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[10][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[10][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[10][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[10][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[10][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[10][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[11][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[11][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[11][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[11][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[11][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[11][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[11][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[11][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[11][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[11][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[11][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[11][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[11][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[11][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[11][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[11][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[11][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[11][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[11][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[11][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[11][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[11][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[11][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[11][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[11][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[11][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[11][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[11][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[11][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[11][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[11][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[11][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[11][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[11][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[11][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[11][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[11][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[11][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[11][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[11][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[11][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[12][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[12][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[12][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[12][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[12][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[12][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[12][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[12][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[12][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[12][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[12][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[12][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[12][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[12][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[12][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[12][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[12][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[12][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[12][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[12][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[12][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[12][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[12][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[12][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[12][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[12][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[12][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[12][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[12][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[12][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[12][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[12][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[12][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[12][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[12][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[12][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[12][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[12][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[12][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[12][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[12][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[13][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[13][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[13][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[13][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[13][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[13][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[13][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[13][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[13][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[13][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[13][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[13][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[13][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[13][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[13][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[13][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[13][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[13][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[13][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[13][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[13][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[13][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[13][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[13][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[13][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[13][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[13][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[13][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[13][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[13][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[13][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[13][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[13][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[13][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[13][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[13][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[13][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[13][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[13][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[13][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[13][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[14][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[14][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[14][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[14][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[14][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[14][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[14][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[14][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[14][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[14][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[14][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[14][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[14][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[14][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[14][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[14][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[14][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[14][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[14][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[14][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[14][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[14][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[14][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[14][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[14][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[14][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[14][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[14][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[14][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[14][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[14][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[14][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[14][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[14][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[14][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[14][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[14][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[14][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[14][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[14][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[14][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[15][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[15][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[15][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[15][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[15][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[15][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[15][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[15][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[15][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[15][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[15][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[15][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[15][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[15][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[15][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[15][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[15][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[15][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[15][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[15][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[15][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[15][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[15][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[15][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[15][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[15][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[15][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[15][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[15][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[15][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[15][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[15][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[15][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[15][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[15][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[15][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[15][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[15][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[15][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[15][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[15][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[16][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[16][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[16][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[16][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[16][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[16][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[16][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[16][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[16][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[16][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[16][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[16][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[16][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[16][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[16][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[16][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[16][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[16][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[16][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[16][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[16][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[16][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[16][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[16][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[16][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[16][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[16][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[16][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[16][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[16][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[16][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[16][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[16][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[16][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[16][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[16][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[16][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[16][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[16][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[16][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[16][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[17][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[17][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[17][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[17][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[17][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[17][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[17][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[17][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[17][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[17][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[17][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[17][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[17][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[17][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[17][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[17][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[17][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[17][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[17][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[17][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[17][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[17][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[17][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[17][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[17][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[17][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[17][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[17][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[17][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[17][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[17][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[17][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[17][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[17][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[17][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[17][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[17][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[17][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[17][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[17][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[17][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[18][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[18][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[18][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[18][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[18][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[18][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[18][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[18][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[18][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[18][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[18][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[18][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[18][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[18][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[18][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[18][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[18][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[18][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[18][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[18][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[18][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[18][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[18][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[18][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[18][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[18][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[18][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[18][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[18][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[18][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[18][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[18][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[18][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[18][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[18][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[18][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[18][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[18][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[18][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[18][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[18][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[19][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[19][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[19][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[19][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[19][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[19][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[19][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[19][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[19][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[19][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[19][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[19][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[19][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[19][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[19][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[19][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[19][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[19][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[19][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[19][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[19][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[19][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[19][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[19][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[19][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[19][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[19][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[19][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[19][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[19][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[19][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[19][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[19][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[19][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[19][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[19][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[19][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[19][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[19][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[19][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[19][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[20][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[20][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[20][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[20][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[20][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[20][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[20][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[20][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[20][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[20][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[20][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[20][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[20][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[20][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[20][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[20][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[20][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[20][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[20][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[20][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[20][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[20][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[20][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[20][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[20][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[20][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[20][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[20][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[20][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[20][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[20][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[20][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[20][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[20][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[20][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[20][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[20][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[20][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[20][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[20][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[20][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[21][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[21][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[21][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[21][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[21][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[21][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[21][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[21][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[21][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[21][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[21][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[21][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[21][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[21][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[21][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[21][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[21][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[21][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[21][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[21][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[21][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[21][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[21][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[21][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[21][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[21][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[21][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[21][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[21][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[21][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[21][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[21][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[21][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[21][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[21][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[21][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[21][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[21][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[21][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[21][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[21][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[22][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[22][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[22][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[22][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[22][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[22][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[22][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[22][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[22][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[22][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[22][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[22][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[22][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[22][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[22][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[22][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[22][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[22][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[22][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[22][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[22][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[22][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[22][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[22][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[22][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[22][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[22][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[22][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[22][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[22][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[22][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[22][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[22][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[22][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[22][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[22][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[22][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[22][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[22][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[22][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[22][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[23][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[23][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[23][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[23][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[23][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[23][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[23][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[23][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[23][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[23][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[23][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[23][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[23][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[23][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[23][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[23][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[23][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[23][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[23][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[23][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[23][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[23][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[23][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[23][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[23][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[23][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[23][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[23][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[23][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[23][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[23][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[23][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[23][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[23][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[23][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[23][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[23][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[23][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[23][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[23][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[23][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[24][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[24][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[24][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[24][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[24][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[24][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[24][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[24][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[24][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[24][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[24][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[24][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[24][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[24][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[24][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[24][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[24][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[24][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[24][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[24][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[24][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[24][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[24][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[24][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[24][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[24][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[24][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[24][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[24][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[24][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[24][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[24][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[24][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[24][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[24][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[24][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[24][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[24][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[24][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[24][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[24][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[25][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[25][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[25][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[25][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[25][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[25][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[25][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[25][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[25][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[25][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[25][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[25][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[25][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[25][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[25][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[25][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[25][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[25][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[25][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[25][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[25][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[25][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[25][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[25][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[25][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[25][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[25][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[25][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[25][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[25][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[25][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[25][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[25][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[25][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[25][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[25][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[25][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[25][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[25][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[25][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[25][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[26][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[26][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[26][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[26][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[26][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[26][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[26][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[26][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[26][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[26][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[26][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[26][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[26][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[26][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[26][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[26][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[26][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[26][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[26][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[26][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[26][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[26][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[26][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[26][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[26][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[26][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[26][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[26][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[26][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[26][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[26][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[26][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[26][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[26][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[26][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[26][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[26][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[26][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[26][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[26][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[26][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[27][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[27][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[27][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[27][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[27][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[27][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[27][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[27][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[27][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[27][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[27][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[27][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[27][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[27][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[27][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[27][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[27][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[27][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[27][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[27][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[27][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[27][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[27][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[27][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[27][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[27][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[27][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[27][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[27][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[27][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[27][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[27][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[27][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[27][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[27][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[27][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[27][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[27][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[27][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[27][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[27][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[28][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[28][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[28][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[28][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[28][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[28][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[28][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[28][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[28][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[28][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[28][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[28][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[28][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[28][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[28][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[28][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[28][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[28][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[28][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[28][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[28][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[28][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[28][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[28][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[28][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[28][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[28][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[28][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[28][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[28][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[28][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[28][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[28][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[28][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[28][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[28][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[28][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[28][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[28][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[28][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[28][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[29][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[29][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[29][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[29][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[29][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[29][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[29][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[29][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[29][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[29][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[29][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[29][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[29][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[29][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[29][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[29][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[29][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[29][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[29][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[29][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[29][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[29][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[29][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[29][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[29][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[29][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[29][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[29][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[29][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[29][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[29][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[29][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[29][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[29][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[29][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[29][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[29][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[29][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[29][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[29][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[29][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[30][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[30][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[30][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[30][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[30][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[30][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[30][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[30][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[30][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[30][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[30][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[30][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[30][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[30][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[30][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[30][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[30][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[30][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[30][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[30][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[30][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[30][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[30][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[30][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[30][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[30][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[30][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[30][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[30][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[30][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[30][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[30][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[30][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[30][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[30][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[30][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[30][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[30][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[30][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[30][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[30][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[31][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[31][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[31][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[31][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[31][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[31][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[31][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[31][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[31][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[31][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[31][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[31][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[31][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[31][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[31][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[31][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[31][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[31][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[31][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[31][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[31][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[31][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[31][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[31][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[31][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[31][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[31][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[31][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[31][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[31][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[31][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[31][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[31][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[31][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[31][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[31][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[31][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[31][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[31][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[31][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[31][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[32][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[32][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[32][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[32][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[32][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[32][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[32][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[32][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[32][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[32][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[32][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[32][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[32][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[32][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[32][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[32][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[32][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[32][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[32][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[32][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[32][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[32][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[32][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[32][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[32][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[32][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[32][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[32][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[32][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[32][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[32][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[32][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[32][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[32][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[32][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[32][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[32][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[32][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[32][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[32][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[32][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[33][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[33][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[33][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[33][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[33][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[33][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[33][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[33][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[33][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[33][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[33][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[33][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[33][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[33][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[33][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[33][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[33][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[33][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[33][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[33][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[33][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[33][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[33][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[33][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[33][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[33][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[33][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[33][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[33][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[33][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[33][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[33][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[33][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[33][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[33][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[33][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[33][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[33][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[33][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[33][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[33][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[34][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[34][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[34][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[34][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[34][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[34][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[34][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[34][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[34][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[34][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[34][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[34][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[34][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[34][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[34][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[34][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[34][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[34][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[34][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[34][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[34][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[34][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[34][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[34][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[34][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[34][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[34][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[34][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[34][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[34][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[34][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[34][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[34][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[34][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[34][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[34][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[34][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[34][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[34][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[34][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[34][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[35][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[35][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[35][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[35][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[35][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[35][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[35][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[35][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[35][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[35][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[35][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[35][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[35][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[35][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[35][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[35][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[35][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[35][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[35][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[35][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[35][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[35][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[35][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[35][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[35][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[35][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[35][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[35][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[35][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[35][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[35][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[35][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[35][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[35][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[35][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[35][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[35][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[35][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[35][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[35][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[35][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[36][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[36][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[36][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[36][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[36][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[36][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[36][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[36][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[36][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[36][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[36][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[36][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[36][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[36][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[36][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[36][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[36][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[36][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[36][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[36][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[36][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[36][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[36][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[36][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[36][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[36][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[36][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[36][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[36][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[36][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[36][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[36][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[36][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[36][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[36][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[36][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[36][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[36][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[36][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[36][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[36][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[37][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[37][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[37][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[37][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[37][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[37][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[37][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[37][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[37][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[37][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[37][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[37][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[37][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[37][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[37][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[37][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[37][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[37][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[37][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[37][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[37][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[37][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[37][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[37][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[37][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[37][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[37][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[37][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[37][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[37][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[37][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[37][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[37][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[37][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[37][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[37][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[37][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[37][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[37][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[37][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[37][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[38][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[38][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[38][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[38][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[38][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[38][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[38][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[38][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[38][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[38][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[38][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[38][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[38][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[38][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[38][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[38][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[38][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[38][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[38][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[38][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[38][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[38][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[38][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[38][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[38][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[38][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[38][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[38][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[38][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[38][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[38][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[38][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[38][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[38][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[38][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[38][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[38][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[38][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[38][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[38][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[38][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[39][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[39][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[39][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[39][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[39][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[39][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[39][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[39][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[39][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[39][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[39][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[39][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[39][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[39][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[39][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[39][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[39][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[39][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[39][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[39][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[39][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[39][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[39][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[39][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[39][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[39][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[39][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[39][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[39][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[39][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[39][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[39][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[39][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[39][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[39][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[39][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[39][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[39][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[39][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[39][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[39][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[40][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[40][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[40][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[40][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[40][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[40][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[40][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[40][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[40][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[40][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[40][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[40][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[40][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[40][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[40][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[40][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[40][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[40][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[40][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[40][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[40][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[40][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[40][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[40][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[40][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[40][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[40][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[40][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[40][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[40][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[40][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[40][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[40][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[40][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[40][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[40][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[40][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[40][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[40][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[40][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[40][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[41][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[41][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[41][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[41][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[41][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[41][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[41][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[41][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[41][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[41][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[41][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[41][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[41][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[41][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[41][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[41][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[41][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[41][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[41][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[41][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[41][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[41][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[41][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[41][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[41][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[41][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[41][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[41][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[41][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[41][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[41][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[41][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[41][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[41][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[41][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[41][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[41][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[41][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[41][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[41][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[41][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[42][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[42][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[42][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[42][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[42][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[42][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[42][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[42][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[42][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[42][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[42][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[42][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[42][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[42][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[42][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[42][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[42][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[42][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[42][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[42][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[42][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[42][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[42][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[42][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[42][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[42][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[42][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[42][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[42][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[42][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[42][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[42][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[42][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[42][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[42][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[42][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[42][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[42][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[42][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[42][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[42][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[43][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[43][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[43][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[43][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[43][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[43][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[43][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[43][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[43][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[43][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[43][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[43][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[43][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[43][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[43][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[43][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[43][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[43][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[43][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[43][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[43][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[43][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[43][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[43][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[43][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[43][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[43][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[43][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[43][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[43][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[43][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[43][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[43][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[43][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[43][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[43][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[43][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[43][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[43][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[43][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[43][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[44][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[44][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[44][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[44][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[44][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[44][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[44][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[44][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[44][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[44][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[44][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[44][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[44][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[44][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[44][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[44][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[44][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[44][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[44][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[44][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[44][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[44][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[44][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[44][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[44][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[44][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[44][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[44][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[44][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[44][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[44][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[44][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[44][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[44][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[44][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[44][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[44][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[44][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[44][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[44][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[44][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[45][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[45][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[45][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[45][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[45][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[45][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[45][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[45][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[45][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[45][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[45][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[45][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[45][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[45][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[45][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[45][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[45][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[45][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[45][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[45][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[45][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[45][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[45][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[45][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[45][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[45][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[45][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[45][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[45][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[45][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[45][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[45][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[45][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[45][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[45][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[45][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[45][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[45][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[45][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[45][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[45][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[46][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[46][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[46][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[46][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[46][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[46][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[46][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[46][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[46][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[46][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[46][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[46][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[46][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[46][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[46][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[46][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[46][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[46][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[46][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[46][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[46][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[46][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[46][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[46][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[46][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[46][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[46][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[46][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[46][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[46][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[46][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[46][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[46][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[46][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[46][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[46][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[46][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[46][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[46][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[46][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[46][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[47][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[47][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[47][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[47][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[47][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[47][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[47][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[47][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[47][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[47][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[47][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[47][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[47][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[47][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[47][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[47][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[47][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[47][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[47][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[47][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[47][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[47][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[47][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[47][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[47][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[47][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[47][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[47][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[47][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[47][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[47][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[47][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[47][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[47][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[47][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[47][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[47][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[47][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[47][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[47][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[47][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[48][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[48][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[48][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[48][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[48][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[48][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[48][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[48][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[48][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[48][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[48][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[48][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[48][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[48][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[48][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[48][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[48][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[48][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[48][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[48][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[48][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[48][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[48][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[48][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[48][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[48][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[48][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[48][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[48][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[48][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[48][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[48][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[48][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[48][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[48][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[48][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[48][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[48][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[48][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[48][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[48][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[49][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[49][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[49][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[49][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[49][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[49][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[49][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[49][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[49][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[49][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[49][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[49][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[49][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[49][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[49][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[49][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[49][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[49][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[49][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[49][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[49][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[49][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[49][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[49][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[49][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[49][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[49][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[49][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[49][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[49][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[49][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[49][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[49][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[49][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[49][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[49][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[49][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[49][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[49][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[49][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[49][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[50][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[50][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[50][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[50][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[50][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[50][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[50][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[50][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[50][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[50][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[50][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[50][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[50][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[50][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[50][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[50][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[50][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[50][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[50][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[50][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[50][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[50][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[50][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[50][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[50][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[50][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[50][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[50][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[50][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[50][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[50][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[50][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[50][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[50][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[50][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[50][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[50][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[50][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[50][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[50][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[50][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[51][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[51][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[51][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[51][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[51][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[51][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[51][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[51][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[51][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[51][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[51][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[51][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[51][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[51][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[51][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[51][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[51][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[51][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[51][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[51][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[51][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[51][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[51][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[51][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[51][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[51][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[51][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[51][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[51][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[51][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[51][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[51][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[51][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[51][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[51][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[51][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[51][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[51][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[51][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[51][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[51][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[52][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[52][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[52][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[52][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[52][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[52][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[52][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[52][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[52][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[52][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[52][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[52][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[52][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[52][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[52][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[52][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[52][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[52][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[52][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[52][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[52][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[52][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[52][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[52][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[52][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[52][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[52][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[52][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[52][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[52][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[52][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[52][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[52][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[52][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[52][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[52][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[52][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[52][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[52][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[52][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[52][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[53][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[53][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[53][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[53][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[53][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[53][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[53][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[53][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[53][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[53][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[53][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[53][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[53][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[53][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[53][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[53][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[53][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[53][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[53][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[53][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[53][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[53][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[53][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[53][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[53][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[53][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[53][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[53][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[53][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[53][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[53][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[53][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[53][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[53][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[53][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[53][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[53][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[53][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[53][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[53][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[53][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[54][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[54][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[54][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[54][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[54][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[54][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[54][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[54][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[54][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[54][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[54][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[54][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[54][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[54][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[54][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[54][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[54][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[54][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[54][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[54][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[54][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[54][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[54][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[54][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[54][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[54][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[54][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[54][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[54][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[54][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[54][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[54][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[54][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[54][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[54][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[54][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[54][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[54][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[54][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[54][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[54][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[55][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[55][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[55][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[55][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[55][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[55][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[55][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[55][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[55][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[55][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[55][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[55][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[55][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[55][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[55][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[55][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[55][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[55][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[55][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[55][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[55][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[55][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[55][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[55][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[55][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[55][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[55][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[55][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[55][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[55][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[55][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[55][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[55][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[55][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[55][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[55][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[55][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[55][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[55][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[55][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[55][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[56][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[56][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[56][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[56][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[56][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[56][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[56][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[56][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[56][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[56][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[56][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[56][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[56][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[56][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[56][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[56][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[56][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[56][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[56][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[56][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[56][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[56][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[56][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[56][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[56][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[56][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[56][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[56][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[56][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[56][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[56][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[56][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[56][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[56][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[56][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[56][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[56][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[56][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[56][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[56][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[56][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[57][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[57][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[57][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[57][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[57][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[57][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[57][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[57][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[57][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[57][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[57][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[57][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[57][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[57][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[57][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[57][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[57][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[57][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[57][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[57][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[57][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[57][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[57][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[57][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[57][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[57][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[57][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[57][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[57][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[57][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[57][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[57][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[57][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[57][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[57][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[57][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[57][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[57][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[57][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[57][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[57][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[58][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[58][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[58][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[58][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[58][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[58][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[58][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[58][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[58][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[58][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[58][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[58][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[58][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[58][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[58][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[58][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[58][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[58][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[58][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[58][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[58][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[58][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[58][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[58][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[58][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[58][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[58][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[58][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[58][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[58][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[58][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[58][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[58][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[58][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[58][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[58][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[58][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[58][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[58][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[58][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[58][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[59][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[59][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[59][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[59][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[59][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[59][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[59][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[59][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[59][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[59][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[59][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[59][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[59][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[59][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[59][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[59][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[59][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[59][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[59][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[59][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[59][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[59][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[59][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[59][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[59][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[59][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[59][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[59][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[59][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[59][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[59][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[59][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[59][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[59][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[59][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[59][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[59][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[59][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[59][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[59][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[59][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[60][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[60][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[60][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[60][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[60][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[60][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[60][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[60][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[60][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[60][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[60][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[60][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[60][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[60][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[60][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[60][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[60][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[60][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[60][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[60][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[60][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[60][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[60][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[60][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[60][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[60][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[60][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[60][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[60][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[60][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[60][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[60][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[60][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[60][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[60][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[60][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[60][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[60][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[60][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[60][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[60][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[61][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[61][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[61][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[61][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[61][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[61][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[61][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[61][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[61][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[61][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[61][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[61][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[61][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[61][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[61][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[61][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[61][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[61][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[61][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[61][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[61][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[61][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[61][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[61][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[61][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[61][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[61][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[61][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[61][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[61][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[61][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[61][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[61][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[61][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[61][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[61][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[61][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[61][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[61][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[61][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[61][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[62][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[62][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[62][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[62][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[62][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[62][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[62][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[62][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[62][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[62][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[62][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[62][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[62][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[62][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[62][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[62][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[62][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[62][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[62][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[62][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[62][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[62][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[62][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[62][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[62][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[62][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[62][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[62][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[62][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[62][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[62][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[62][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[62][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[62][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[62][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[62][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[62][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[62][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[62][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[62][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[62][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[63][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[63][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[63][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[63][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[63][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[63][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[63][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[63][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[63][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[63][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[63][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[63][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[63][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[63][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[63][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[63][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[63][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[63][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[63][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[63][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[63][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[63][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[63][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[63][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[63][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[63][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[63][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[63][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[63][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[63][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[63][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[63][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[63][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[63][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[63][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[63][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[63][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[63][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[63][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[63][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[63][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[64][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[64][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[64][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[64][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[64][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[64][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[64][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[64][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[64][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[64][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[64][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[64][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[64][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[64][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[64][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[64][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[64][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[64][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[64][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[64][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[64][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[64][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[64][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[64][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[64][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[64][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[64][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[64][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[64][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[64][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[64][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[64][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[64][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[64][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[64][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[64][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[64][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[64][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[64][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[64][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[64][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[65][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[65][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[65][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[65][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[65][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[65][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[65][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[65][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[65][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[65][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[65][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[65][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[65][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[65][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[65][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[65][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[65][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[65][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[65][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[65][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[65][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[65][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[65][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[65][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[65][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[65][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[65][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[65][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[65][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[65][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[65][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[65][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[65][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[65][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[65][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[65][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[65][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[65][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[65][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[65][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[65][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[66][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[66][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[66][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[66][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[66][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[66][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[66][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[66][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[66][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[66][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[66][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[66][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[66][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[66][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[66][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[66][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[66][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[66][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[66][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[66][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[66][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[66][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[66][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[66][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[66][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[66][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[66][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[66][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[66][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[66][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[66][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[66][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[66][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[66][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[66][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[66][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[66][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[66][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[66][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[66][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[66][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[67][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[67][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[67][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[67][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[67][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[67][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[67][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[67][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[67][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[67][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[67][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[67][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[67][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[67][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[67][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[67][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[67][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[67][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[67][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[67][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[67][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[67][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[67][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[67][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[67][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[67][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[67][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[67][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[67][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[67][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[67][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[67][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[67][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[67][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[67][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[67][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[67][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[67][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[67][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[67][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[67][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[68][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[68][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[68][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[68][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[68][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[68][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[68][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[68][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[68][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[68][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[68][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[68][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[68][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[68][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[68][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[68][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[68][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[68][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[68][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[68][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[68][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[68][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[68][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[68][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[68][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[68][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[68][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[68][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[68][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[68][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[68][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[68][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[68][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[68][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[68][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[68][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[68][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[68][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[68][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[68][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[68][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[69][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[69][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[69][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[69][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[69][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[69][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[69][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[69][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[69][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[69][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[69][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[69][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[69][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[69][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[69][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[69][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[69][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[69][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[69][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[69][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[69][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[69][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[69][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[69][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[69][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[69][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[69][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[69][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[69][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[69][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[69][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[69][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[69][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[69][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[69][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[69][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[69][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[69][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[69][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[69][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[69][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[70][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[70][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[70][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[70][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[70][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[70][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[70][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[70][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[70][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[70][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[70][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[70][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[70][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[70][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[70][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[70][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[70][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[70][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[70][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[70][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[70][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[70][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[70][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[70][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[70][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[70][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[70][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[70][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[70][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[70][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[70][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[70][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[70][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[70][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[70][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[70][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[70][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[70][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[70][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[70][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[70][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[71][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[71][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[71][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[71][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[71][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[71][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[71][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[71][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[71][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[71][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[71][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[71][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[71][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[71][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[71][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[71][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[71][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[71][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[71][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[71][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[71][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[71][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[71][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[71][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[71][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[71][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[71][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[71][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[71][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[71][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[71][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[71][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[71][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[71][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[71][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[71][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[71][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[71][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[71][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[71][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[71][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[72][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[72][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[72][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[72][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[72][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[72][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[72][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[72][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[72][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[72][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[72][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[72][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[72][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[72][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[72][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[72][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[72][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[72][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[72][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[72][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[72][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[72][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[72][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[72][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[72][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[72][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[72][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[72][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[72][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[72][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[72][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[72][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[72][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[72][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[72][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[72][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[72][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[72][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[72][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[72][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[72][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[73][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[73][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[73][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[73][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[73][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[73][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[73][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[73][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[73][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[73][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[73][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[73][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[73][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[73][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[73][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[73][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[73][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[73][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[73][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[73][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[73][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[73][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[73][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[73][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[73][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[73][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[73][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[73][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[73][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[73][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[73][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[73][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[73][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[73][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[73][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[73][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[73][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[73][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[73][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[73][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[73][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[74][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[74][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[74][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[74][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[74][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[74][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[74][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[74][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[74][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[74][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[74][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[74][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[74][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[74][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[74][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[74][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[74][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[74][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[74][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[74][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[74][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[74][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[74][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[74][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[74][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[74][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[74][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[74][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[74][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[74][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[74][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[74][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[74][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[74][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[74][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[74][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[74][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[74][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[74][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[74][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[74][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[75][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[75][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[75][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[75][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[75][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[75][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[75][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[75][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[75][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[75][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[75][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[75][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[75][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[75][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[75][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[75][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[75][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[75][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[75][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[75][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[75][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[75][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[75][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[75][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[75][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[75][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[75][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[75][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[75][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[75][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[75][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[75][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[75][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[75][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[75][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[75][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[75][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[75][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[75][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[75][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[75][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[76][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[76][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[76][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[76][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[76][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[76][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[76][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[76][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[76][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[76][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[76][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[76][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[76][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[76][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[76][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[76][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[76][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[76][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[76][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[76][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[76][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[76][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[76][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[76][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[76][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[76][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[76][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[76][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[76][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[76][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[76][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[76][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[76][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[76][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[76][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[76][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[76][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[76][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[76][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[76][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[76][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[77][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[77][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[77][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[77][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[77][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[77][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[77][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[77][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[77][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[77][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[77][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[77][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[77][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[77][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[77][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[77][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[77][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[77][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[77][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[77][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[77][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[77][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[77][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[77][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[77][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[77][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[77][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[77][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[77][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[77][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[77][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[77][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[77][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[77][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[77][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[77][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[77][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[77][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[77][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[77][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[77][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[78][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[78][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[78][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[78][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[78][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[78][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[78][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[78][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[78][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[78][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[78][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[78][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[78][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[78][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[78][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[78][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[78][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[78][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[78][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[78][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[78][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[78][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[78][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[78][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[78][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[78][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[78][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[78][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[78][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[78][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[78][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[78][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[78][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[78][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[78][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[78][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[78][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[78][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[78][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[78][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[78][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[79][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[79][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[79][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[79][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[79][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[79][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[79][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[79][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[79][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[79][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[79][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[79][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[79][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[79][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[79][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[79][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[79][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[79][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[79][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[79][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[79][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[79][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[79][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[79][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[79][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[79][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[79][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[79][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[79][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[79][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[79][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[79][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[79][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[79][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[79][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[79][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[79][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[79][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[79][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[79][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[79][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[80][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[80][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[80][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[80][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[80][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[80][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[80][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[80][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[80][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[80][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[80][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[80][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[80][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[80][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[80][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[80][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[80][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[80][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[80][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[80][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[80][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[80][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[80][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[80][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[80][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[80][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[80][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[80][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[80][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[80][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[80][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[80][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[80][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[80][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[80][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[80][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[80][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[80][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[80][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[80][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[80][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[81][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[81][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[81][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[81][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[81][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[81][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[81][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[81][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[81][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[81][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[81][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[81][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[81][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[81][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[81][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[81][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[81][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[81][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[81][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[81][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[81][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[81][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[81][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[81][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[81][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[81][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[81][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[81][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[81][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[81][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[81][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[81][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[81][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[81][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[81][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[81][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[81][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[81][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[81][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[81][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[81][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[82][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[82][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[82][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[82][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[82][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[82][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[82][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[82][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[82][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[82][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[82][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[82][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[82][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[82][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[82][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[82][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[82][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[82][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[82][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[82][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[82][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[82][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[82][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[82][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[82][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[82][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[82][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[82][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[82][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[82][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[82][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[82][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[82][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[82][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[82][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[82][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[82][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[82][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[82][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[82][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[82][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[83][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[83][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[83][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[83][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[83][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[83][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[83][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[83][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[83][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[83][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[83][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[83][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[83][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[83][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[83][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[83][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[83][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[83][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[83][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[83][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[83][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[83][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[83][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[83][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[83][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[83][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[83][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[83][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[83][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[83][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[83][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[83][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[83][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[83][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[83][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[83][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[83][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[83][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[83][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[83][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[83][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[84][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[84][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[84][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[84][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[84][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[84][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[84][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[84][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[84][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[84][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[84][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[84][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[84][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[84][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[84][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[84][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[84][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[84][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[84][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[84][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[84][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[84][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[84][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[84][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[84][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[84][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[84][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[84][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[84][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[84][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[84][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[84][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[84][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[84][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[84][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[84][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[84][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[84][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[84][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[84][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[84][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[85][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[85][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[85][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[85][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[85][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[85][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[85][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[85][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[85][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[85][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[85][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[85][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[85][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[85][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[85][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[85][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[85][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[85][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[85][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[85][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[85][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[85][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[85][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[85][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[85][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[85][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[85][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[85][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[85][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[85][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[85][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[85][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[85][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[85][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[85][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[85][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[85][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[85][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[85][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[85][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[85][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[86][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[86][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[86][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[86][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[86][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[86][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[86][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[86][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[86][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[86][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[86][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[86][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[86][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[86][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[86][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[86][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[86][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[86][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[86][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[86][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[86][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[86][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[86][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[86][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[86][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[86][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[86][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[86][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[86][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[86][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[86][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[86][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[86][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[86][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[86][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[86][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[86][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[86][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[86][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[86][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[86][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[87][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[87][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[87][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[87][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[87][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[87][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[87][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[87][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[87][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[87][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[87][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[87][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[87][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[87][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[87][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[87][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[87][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[87][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[87][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[87][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[87][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[87][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[87][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[87][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[87][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[87][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[87][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[87][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[87][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[87][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[87][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[87][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[87][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[87][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[87][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[87][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[87][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[87][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[87][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[87][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[87][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[88][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[88][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[88][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[88][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[88][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[88][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[88][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[88][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[88][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[88][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[88][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[88][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[88][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[88][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[88][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[88][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[88][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[88][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[88][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[88][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[88][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[88][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[88][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[88][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[88][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[88][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[88][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[88][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[88][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[88][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[88][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[88][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[88][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[88][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[88][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[88][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[88][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[88][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[88][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[88][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[88][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[89][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[89][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[89][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[89][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[89][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[89][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[89][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[89][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[89][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[89][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[89][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[89][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[89][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[89][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[89][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[89][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[89][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[89][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[89][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[89][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[89][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[89][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[89][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[89][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[89][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[89][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[89][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[89][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[89][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[89][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[89][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[89][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[89][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[89][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[89][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[89][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[89][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[89][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[89][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[89][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[89][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[90][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[90][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[90][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[90][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[90][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[90][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[90][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[90][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[90][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[90][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[90][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[90][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[90][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[90][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[90][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[90][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[90][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[90][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[90][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[90][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[90][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[90][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[90][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[90][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[90][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[90][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[90][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[90][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[90][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[90][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[90][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[90][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[90][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[90][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[90][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[90][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[90][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[90][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[90][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[90][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[90][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[91][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[91][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[91][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[91][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[91][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[91][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[91][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[91][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[91][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[91][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[91][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[91][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[91][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[91][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[91][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[91][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[91][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[91][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[91][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[91][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[91][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[91][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[91][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[91][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[91][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[91][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[91][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[91][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[91][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[91][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[91][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[91][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[91][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[91][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[91][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[91][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[91][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[91][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[91][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[91][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[91][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[92][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[92][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[92][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[92][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[92][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[92][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[92][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[92][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[92][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[92][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[92][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[92][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[92][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[92][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[92][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[92][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[92][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[92][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[92][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[92][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[92][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[92][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[92][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[92][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[92][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[92][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[92][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[92][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[92][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[92][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[92][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[92][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[92][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[92][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[92][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[92][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[92][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[92][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[92][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[92][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[92][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[93][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[93][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[93][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[93][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[93][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[93][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[93][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[93][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[93][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[93][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[93][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[93][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[93][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[93][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[93][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[93][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[93][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[93][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[93][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[93][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[93][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[93][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[93][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[93][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[93][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[93][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[93][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[93][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[93][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[93][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[93][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[93][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[93][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[93][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[93][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[93][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[93][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[93][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[93][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[93][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[93][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[94][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[94][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[94][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[94][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[94][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[94][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[94][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[94][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[94][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[94][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[94][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[94][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[94][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[94][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[94][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[94][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[94][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[94][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[94][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[94][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[94][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[94][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[94][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[94][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[94][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[94][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[94][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[94][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[94][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[94][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[94][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[94][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[94][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[94][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[94][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[94][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[94][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[94][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[94][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[94][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[94][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[95][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[95][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[95][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[95][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[95][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[95][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[95][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[95][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[95][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[95][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[95][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[95][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[95][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[95][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[95][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[95][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[95][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[95][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[95][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[95][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[95][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[95][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[95][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[95][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[95][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[95][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[95][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[95][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[95][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[95][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[95][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[95][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[95][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[95][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[95][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[95][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[95][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[95][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[95][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[95][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[95][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[96][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[96][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[96][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[96][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[96][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[96][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[96][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[96][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[96][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[96][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[96][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[96][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[96][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[96][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[96][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[96][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[96][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[96][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[96][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[96][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[96][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[96][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[96][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[96][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[96][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[96][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[96][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[96][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[96][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[96][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[96][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[96][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[96][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[96][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[96][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[96][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[96][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[96][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[96][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[96][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[96][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[97][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[97][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[97][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[97][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[97][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[97][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[97][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[97][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[97][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[97][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[97][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[97][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[97][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[97][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[97][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[97][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[97][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[97][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[97][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[97][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[97][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[97][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[97][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[97][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[97][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[97][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[97][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[97][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[97][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[97][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[97][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[97][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[97][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[97][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[97][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[97][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[97][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[97][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[97][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[97][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[97][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[98][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[98][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[98][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[98][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[98][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[98][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[98][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[98][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[98][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[98][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[98][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[98][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[98][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[98][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[98][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[98][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[98][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[98][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[98][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[98][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[98][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[98][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[98][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[98][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[98][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[98][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[98][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[98][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[98][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[98][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[98][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[98][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[98][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[98][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[98][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[98][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[98][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[98][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[98][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[98][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[98][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[99][0]~FF  (.D(\data_to_tx_packet_reg[0] ), .CE(\i15/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[99][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[99][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[99][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[99][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[99][1]~FF  (.D(\data_to_tx_packet_reg[1] ), .CE(\i15/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[99][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[99][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[99][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[99][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[99][2]~FF  (.D(\data_to_tx_packet_reg[2] ), .CE(\i15/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[99][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[99][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[99][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[99][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[99][3]~FF  (.D(\data_to_tx_packet_reg[3] ), .CE(\i15/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[99][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[99][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[99][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[99][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[99][4]~FF  (.D(\data_to_tx_packet_reg[4] ), .CE(\i15/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[99][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[99][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[99][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[99][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[99][5]~FF  (.D(\data_to_tx_packet_reg[5] ), .CE(\i15/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[99][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[99][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[99][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[99][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[99][6]~FF  (.D(\data_to_tx_packet_reg[6] ), .CE(\i15/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[99][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[99][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[99][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[99][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[99][7]~FF  (.D(\data_to_tx_packet_reg[7] ), .CE(\i15/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[99][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[99][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[99][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[99][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[99][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[100][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[100][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[100][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[100][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[100][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[100][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[100][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[100][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[100][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[100][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[100][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[100][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[100][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[100][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[100][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[100][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[100][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[100][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[100][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[100][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[100][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[100][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[100][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[100][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[100][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[100][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[100][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[100][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[100][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[100][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[100][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[100][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[100][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[100][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[100][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[100][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[100][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[100][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[100][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[100][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[100][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[101][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[101][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[101][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[101][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[101][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[101][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[101][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[101][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[101][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[101][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[101][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[101][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[101][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[101][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[101][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[101][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[101][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[101][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[101][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[101][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[101][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[101][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[101][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[101][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[101][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[101][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[101][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[101][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[101][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[101][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[101][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[101][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[101][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[101][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[101][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[101][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[101][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[101][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[101][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[101][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[101][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[102][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[102][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[102][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[102][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[102][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[102][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[102][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[102][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[102][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[102][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[102][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[102][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[102][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[102][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[102][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[102][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[102][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[102][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[102][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[102][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[102][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[102][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[102][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[102][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[102][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[102][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[102][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[102][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[102][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[102][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[102][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[102][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[102][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[102][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[102][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[102][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[102][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[102][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[102][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[102][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[102][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[103][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[103][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[103][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[103][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[103][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[103][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[103][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[103][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[103][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[103][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[103][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[103][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[103][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[103][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[103][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[103][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[103][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[103][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[103][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[103][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[103][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[103][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[103][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[103][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[103][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[103][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[103][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[103][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[103][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[103][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[103][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[103][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[103][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[103][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[103][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[103][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[103][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[103][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[103][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[103][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[103][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[104][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[104][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[104][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[104][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[104][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[104][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[104][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[104][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[104][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[104][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[104][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[104][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[104][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[104][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[104][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[104][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[104][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[104][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[104][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[104][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[104][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[104][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[104][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[104][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[104][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[104][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[104][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[104][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[104][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[104][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[104][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[104][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[104][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[104][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[104][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[104][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[104][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[104][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[104][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[104][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[104][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[105][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[105][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[105][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[105][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[105][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[105][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[105][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[105][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[105][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[105][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[105][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[105][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[105][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[105][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[105][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[105][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[105][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[105][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[105][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[105][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[105][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[105][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[105][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[105][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[105][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[105][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[105][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[105][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[105][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[105][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[105][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[105][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[105][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[105][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[105][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[105][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[105][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[105][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[105][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[105][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[105][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[106][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[106][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[106][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[106][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[106][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[106][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[106][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[106][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[106][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[106][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[106][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[106][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[106][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[106][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[106][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[106][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[106][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[106][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[106][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[106][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[106][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[106][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[106][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[106][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[106][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[106][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[106][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[106][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[106][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[106][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[106][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[106][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[106][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[106][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[106][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[106][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[106][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[106][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[106][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[106][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[106][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[107][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[107][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[107][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[107][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[107][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[107][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[107][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[107][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[107][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[107][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[107][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[107][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[107][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[107][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[107][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[107][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[107][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[107][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[107][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[107][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[107][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[107][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[107][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[107][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[107][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[107][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[107][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[107][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[107][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[107][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[107][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[107][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[107][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[107][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[107][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[107][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[107][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[107][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[107][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[107][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[107][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[108][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[108][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[108][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[108][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[108][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[108][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[108][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[108][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[108][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[108][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[108][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[108][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[108][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[108][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[108][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[108][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[108][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[108][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[108][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[108][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[108][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[108][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[108][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[108][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[108][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[108][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[108][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[108][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[108][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[108][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[108][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[108][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[108][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[108][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[108][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[108][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[108][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[108][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[108][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[108][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[108][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[109][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[109][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[109][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[109][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[109][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[109][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[109][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[109][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[109][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[109][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[109][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[109][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[109][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[109][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[109][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[109][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[109][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[109][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[109][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[109][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[109][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[109][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[109][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[109][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[109][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[109][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[109][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[109][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[109][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[109][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[109][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[109][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[109][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[109][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[109][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[109][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[109][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[109][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[109][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[109][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[109][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[110][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[110][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[110][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[110][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[110][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[110][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[110][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[110][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[110][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[110][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[110][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[110][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[110][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[110][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[110][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[110][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[110][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[110][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[110][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[110][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[110][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[110][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[110][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[110][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[110][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[110][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[110][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[110][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[110][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[110][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[110][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[110][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[110][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[110][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[110][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[110][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[110][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[110][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[110][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[110][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[110][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[111][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[111][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[111][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[111][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[111][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[111][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[111][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[111][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[111][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[111][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[111][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[111][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[111][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[111][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[111][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[111][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[111][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[111][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[111][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[111][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[111][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[111][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[111][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[111][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[111][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[111][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[111][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[111][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[111][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[111][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[111][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[111][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[111][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[111][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[111][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[111][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[111][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[111][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[111][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[111][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[111][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[112][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[112][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[112][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[112][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[112][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[112][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[112][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[112][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[112][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[112][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[112][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[112][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[112][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[112][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[112][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[112][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[112][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[112][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[112][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[112][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[112][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[112][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[112][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[112][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[112][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[112][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[112][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[112][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[112][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[112][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[112][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[112][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[112][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[112][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[112][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[112][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[112][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[112][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[112][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[112][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[112][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[113][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[113][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[113][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[113][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[113][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[113][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[113][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[113][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[113][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[113][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[113][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[113][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[113][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[113][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[113][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[113][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[113][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[113][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[113][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[113][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[113][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[113][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[113][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[113][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[113][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[113][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[113][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[113][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[113][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[113][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[113][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[113][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[113][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[113][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[113][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[113][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[113][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[113][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[113][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[113][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[113][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[114][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[114][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[114][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[114][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[114][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[114][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[114][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[114][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[114][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[114][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[114][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[114][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[114][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[114][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[114][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[114][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[114][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[114][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[114][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[114][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[114][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[114][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[114][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[114][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[114][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[114][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[114][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[114][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[114][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[114][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[114][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[114][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[114][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[114][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[114][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[114][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[114][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[114][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[114][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[114][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[114][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[115][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[115][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[115][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[115][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[115][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[115][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[115][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[115][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[115][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[115][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[115][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[115][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[115][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[115][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[115][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[115][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[115][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[115][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[115][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[115][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[115][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[115][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[115][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[115][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[115][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[115][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[115][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[115][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[115][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[115][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[115][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[115][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[115][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[115][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[115][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[115][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[115][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[115][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[115][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[115][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[115][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[116][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[116][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[116][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[116][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[116][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[116][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[116][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[116][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[116][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[116][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[116][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[116][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[116][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[116][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[116][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[116][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[116][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[116][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[116][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[116][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[116][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[116][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[116][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[116][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[116][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[116][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[116][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[116][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[116][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[116][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[116][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[116][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[116][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[116][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[116][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[116][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[116][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[116][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[116][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[116][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[116][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[117][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[117][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[117][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[117][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[117][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[117][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[117][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[117][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[117][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[117][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[117][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[117][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[117][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[117][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[117][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[117][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[117][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[117][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[117][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[117][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[117][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[117][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[117][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[117][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[117][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[117][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[117][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[117][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[117][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[117][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[117][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[117][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[117][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[117][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[117][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[117][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[117][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[117][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[117][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[117][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[117][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[118][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[118][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[118][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[118][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[118][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[118][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[118][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[118][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[118][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[118][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[118][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[118][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[118][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[118][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[118][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[118][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[118][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[118][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[118][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[118][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[118][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[118][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[118][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[118][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[118][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[118][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[118][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[118][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[118][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[118][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[118][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[118][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[118][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[118][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[118][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[118][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[118][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[118][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[118][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[118][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[118][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[119][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[119][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[119][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[119][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[119][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[119][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[119][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[119][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[119][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[119][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[119][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[119][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[119][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[119][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[119][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[119][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[119][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[119][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[119][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[119][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[119][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[119][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[119][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[119][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[119][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[119][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[119][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[119][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[119][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[119][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[119][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[119][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[119][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[119][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[119][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[119][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[119][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[119][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[119][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[119][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[119][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[120][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[120][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[120][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[120][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[120][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[120][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[120][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[120][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[120][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[120][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[120][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[120][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[120][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[120][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[120][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[120][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[120][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[120][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[120][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[120][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[120][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[120][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[120][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[120][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[120][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[120][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[120][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[120][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[120][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[120][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[120][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[120][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[120][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[120][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[120][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[120][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[120][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[120][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[120][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[120][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[120][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[121][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[121][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[121][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[121][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[121][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[121][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[121][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[121][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[121][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[121][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[121][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[121][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[121][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[121][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[121][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[121][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[121][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[121][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[121][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[121][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[121][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[121][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[121][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[121][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[121][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[121][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[121][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[121][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[121][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[121][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[121][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[121][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[121][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[121][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[121][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[121][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[121][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[121][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[121][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[121][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[121][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[122][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[122][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[122][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[122][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[122][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[122][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[122][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[122][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[122][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[122][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[122][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[122][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[122][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[122][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[122][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[122][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[122][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[122][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[122][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[122][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[122][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[122][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[122][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[122][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[122][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[122][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[122][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[122][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[122][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[122][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[122][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[122][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[122][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[122][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[122][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[122][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[122][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[122][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[122][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[122][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[122][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[123][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[123][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[123][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[123][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[123][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[123][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[123][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[123][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[123][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[123][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[123][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[123][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[123][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[123][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[123][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[123][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[123][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[123][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[123][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[123][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[123][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[123][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[123][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[123][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[123][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[123][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[123][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[123][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[123][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[123][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[123][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[123][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[123][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[123][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[123][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[123][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[123][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[123][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[123][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[123][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[123][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[124][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[124][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[124][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[124][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[124][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[124][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[124][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[124][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[124][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[124][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[124][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[124][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[124][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[124][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[124][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[124][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[124][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[124][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[124][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[124][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[124][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[124][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[124][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[124][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[124][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[124][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[124][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[124][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[124][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[124][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[124][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[124][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[124][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[124][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[124][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[124][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[124][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[124][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[124][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[124][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[124][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[125][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[125][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[125][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[125][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[125][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[125][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[125][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[125][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[125][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[125][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[125][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[125][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[125][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[125][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[125][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[125][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[125][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[125][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[125][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[125][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[125][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[125][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[125][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[125][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[125][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[125][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[125][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[125][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[125][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[125][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[125][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[125][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[125][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[125][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[125][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[125][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[125][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[125][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[125][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[125][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[125][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[126][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[126][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[126][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[126][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[126][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[126][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[126][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[126][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[126][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[126][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[126][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[126][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[126][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[126][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[126][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[126][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[126][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[126][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[126][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[126][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[126][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[126][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[126][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[126][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[126][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[126][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[126][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[126][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[126][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[126][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[126][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[126][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[126][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[126][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[126][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[126][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[126][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[126][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[126][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[126][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[126][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[127][0]~FF  (.D(\data_to_tx_packet_reg[0] ), 
           .CE(\i15/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[127][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[127][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][0]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][0]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][0]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][0]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[127][0]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[127][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[127][1]~FF  (.D(\data_to_tx_packet_reg[1] ), 
           .CE(\i15/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[127][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[127][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][1]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][1]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][1]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][1]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[127][1]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[127][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[127][2]~FF  (.D(\data_to_tx_packet_reg[2] ), 
           .CE(\i15/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[127][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[127][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][2]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][2]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][2]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][2]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[127][2]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[127][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[127][3]~FF  (.D(\data_to_tx_packet_reg[3] ), 
           .CE(\i15/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[127][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[127][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][3]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][3]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][3]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][3]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[127][3]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[127][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[127][4]~FF  (.D(\data_to_tx_packet_reg[4] ), 
           .CE(\i15/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[127][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[127][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][4]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][4]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][4]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][4]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[127][4]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[127][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[127][5]~FF  (.D(\data_to_tx_packet_reg[5] ), 
           .CE(\i15/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[127][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[127][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][5]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][5]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][5]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][5]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[127][5]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[127][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[127][6]~FF  (.D(\data_to_tx_packet_reg[6] ), 
           .CE(\i15/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[127][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[127][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][6]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][6]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][6]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][6]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[127][6]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[127][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i15/tx_fifo/buff[127][7]~FF  (.D(\data_to_tx_packet_reg[7] ), 
           .CE(\i15/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i15/tx_fifo/buff[127][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i15/tx_fifo/buff[127][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][7]~FF .CE_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][7]~FF .SR_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][7]~FF .D_POLARITY = 1'b1;
    defparam \i15/tx_fifo/buff[127][7]~FF .SR_SYNC = 1'b1;
    defparam \i15/tx_fifo/buff[127][7]~FF .SR_VALUE = 1'b0;
    defparam \i15/tx_fifo/buff[127][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[0][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[0][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[0][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[0][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[0][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[0][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[0][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[0][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[0][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[0][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[0][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[0][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[0][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[0][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[0][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n132 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[0][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[0][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[1][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[1][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[1][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[1][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[1][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[1][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[1][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[1][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[1][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[1][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[1][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[1][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[1][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[1][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[1][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[1][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[1][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[1][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[1][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[1][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[1][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[1][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[1][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[1][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[1][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[1][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[1][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[1][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[1][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[1][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[1][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[1][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[1][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[1][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[1][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[1][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n131 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[1][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[1][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[1][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[1][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[1][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[2][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[2][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[2][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[2][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[2][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[2][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[2][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[2][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[2][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[2][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[2][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[2][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[2][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[2][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[2][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[2][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[2][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[2][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[2][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[2][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[2][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[2][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[2][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[2][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[2][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[2][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[2][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[2][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[2][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[2][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[2][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[2][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[2][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[2][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[2][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[2][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n130 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[2][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[2][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[2][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[2][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[2][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[3][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[3][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[3][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[3][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[3][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[3][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[3][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[3][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[3][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[3][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[3][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[3][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[3][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[3][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[3][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[3][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[3][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[3][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[3][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[3][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[3][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[3][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[3][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[3][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[3][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[3][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[3][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[3][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[3][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[3][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[3][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[3][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[3][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[3][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[3][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[3][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n129 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[3][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[3][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[3][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[3][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[3][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[4][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[4][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[4][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[4][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[4][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[4][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[4][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[4][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[4][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[4][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[4][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[4][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[4][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[4][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[4][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[4][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[4][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[4][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[4][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[4][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[4][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[4][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[4][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[4][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[4][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[4][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[4][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[4][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[4][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[4][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[4][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[4][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[4][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[4][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[4][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[4][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n128 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[4][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[4][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[4][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[4][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[4][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[5][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[5][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[5][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[5][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[5][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[5][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[5][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[5][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[5][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[5][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[5][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[5][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[5][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[5][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[5][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[5][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[5][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[5][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[5][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[5][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[5][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[5][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[5][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[5][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[5][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[5][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[5][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[5][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[5][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[5][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[5][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[5][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[5][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[5][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[5][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[5][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n127 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[5][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[5][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[5][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[5][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[5][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[6][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[6][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[6][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[6][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[6][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[6][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[6][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[6][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[6][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[6][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[6][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[6][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[6][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[6][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[6][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[6][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[6][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[6][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[6][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[6][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[6][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[6][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[6][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[6][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[6][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[6][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[6][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[6][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[6][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[6][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[6][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[6][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[6][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[6][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[6][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[6][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n126 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[6][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[6][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[6][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[6][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[6][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[7][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[7][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[7][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[7][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[7][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[7][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[7][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[7][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[7][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[7][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[7][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[7][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[7][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[7][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[7][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[7][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[7][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[7][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[7][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[7][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[7][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[7][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[7][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[7][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[7][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[7][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[7][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[7][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[7][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[7][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[7][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[7][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[7][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[7][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[7][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[7][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n125 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[7][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[7][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[7][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[7][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[7][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[8][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[8][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[8][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[8][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[8][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[8][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[8][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[8][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[8][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[8][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[8][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[8][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[8][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[8][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[8][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[8][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[8][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[8][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[8][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[8][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[8][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[8][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[8][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[8][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[8][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[8][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[8][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[8][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[8][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[8][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[8][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[8][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[8][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[8][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[8][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[8][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n124 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[8][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[8][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[8][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[8][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[8][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[9][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[9][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[9][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[9][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[9][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[9][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[9][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[9][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[9][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[9][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[9][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[9][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[9][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[9][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[9][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[9][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[9][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[9][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[9][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[9][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[9][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[9][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[9][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[9][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[9][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[9][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[9][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[9][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[9][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[9][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[9][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[9][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[9][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[9][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[9][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[9][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n123 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[9][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[9][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[9][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[9][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[9][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[10][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[10][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[10][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[10][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[10][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[10][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[10][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[10][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[10][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[10][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[10][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[10][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[10][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[10][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[10][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[10][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[10][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[10][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[10][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[10][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[10][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[10][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[10][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[10][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[10][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[10][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[10][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[10][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[10][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[10][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[10][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[10][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[10][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[10][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[10][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[10][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n122 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[10][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[10][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[10][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[10][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[10][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[11][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[11][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[11][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[11][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[11][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[11][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[11][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[11][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[11][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[11][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[11][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[11][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[11][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[11][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[11][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[11][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[11][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[11][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[11][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[11][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[11][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[11][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[11][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[11][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[11][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[11][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[11][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[11][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[11][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[11][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[11][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[11][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[11][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[11][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[11][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[11][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n121 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[11][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[11][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[11][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[11][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[11][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[12][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[12][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[12][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[12][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[12][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[12][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[12][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[12][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[12][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[12][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[12][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[12][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[12][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[12][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[12][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[12][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[12][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[12][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[12][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[12][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[12][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[12][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[12][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[12][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[12][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[12][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[12][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[12][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[12][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[12][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[12][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[12][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[12][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[12][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[12][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[12][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n120 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[12][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[12][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[12][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[12][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[12][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[13][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[13][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[13][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[13][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[13][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[13][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[13][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[13][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[13][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[13][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[13][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[13][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[13][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[13][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[13][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[13][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[13][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[13][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[13][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[13][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[13][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[13][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[13][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[13][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[13][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[13][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[13][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[13][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[13][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[13][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[13][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[13][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[13][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[13][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[13][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[13][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n119 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[13][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[13][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[13][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[13][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[13][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[14][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[14][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[14][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[14][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[14][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[14][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[14][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[14][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[14][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[14][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[14][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[14][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[14][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[14][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[14][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[14][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[14][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[14][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[14][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[14][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[14][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[14][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[14][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[14][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[14][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[14][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[14][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[14][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[14][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[14][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[14][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[14][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[14][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[14][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[14][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[14][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n118 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[14][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[14][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[14][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[14][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[14][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[15][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[15][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[15][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[15][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[15][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[15][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[15][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[15][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[15][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[15][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[15][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[15][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[15][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[15][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[15][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[15][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[15][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[15][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[15][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[15][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[15][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[15][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[15][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[15][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[15][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[15][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[15][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[15][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[15][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[15][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[15][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[15][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[15][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[15][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[15][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[15][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n117 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[15][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[15][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[15][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[15][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[15][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[16][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[16][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[16][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[16][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[16][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[16][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[16][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[16][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[16][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[16][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[16][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[16][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[16][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[16][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[16][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[16][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[16][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[16][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[16][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[16][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[16][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[16][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[16][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[16][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[16][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[16][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[16][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[16][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[16][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[16][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[16][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[16][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[16][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[16][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[16][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[16][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n116 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[16][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[16][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[16][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[16][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[16][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[17][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[17][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[17][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[17][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[17][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[17][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[17][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[17][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[17][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[17][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[17][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[17][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[17][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[17][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[17][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[17][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[17][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[17][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[17][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[17][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[17][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[17][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[17][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[17][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[17][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[17][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[17][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[17][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[17][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[17][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[17][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[17][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[17][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[17][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[17][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[17][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n115 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[17][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[17][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[17][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[17][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[17][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[18][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[18][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[18][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[18][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[18][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[18][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[18][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[18][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[18][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[18][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[18][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[18][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[18][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[18][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[18][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[18][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[18][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[18][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[18][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[18][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[18][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[18][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[18][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[18][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[18][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[18][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[18][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[18][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[18][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[18][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[18][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[18][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[18][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[18][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[18][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[18][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n114 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[18][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[18][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[18][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[18][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[18][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[19][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[19][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[19][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[19][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[19][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[19][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[19][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[19][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[19][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[19][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[19][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[19][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[19][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[19][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[19][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[19][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[19][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[19][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[19][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[19][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[19][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[19][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[19][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[19][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[19][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[19][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[19][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[19][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[19][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[19][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[19][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[19][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[19][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[19][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[19][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[19][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n113 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[19][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[19][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[19][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[19][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[19][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[20][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[20][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[20][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[20][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[20][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[20][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[20][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[20][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[20][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[20][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[20][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[20][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[20][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[20][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[20][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[20][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[20][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[20][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[20][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[20][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[20][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[20][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[20][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[20][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[20][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[20][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[20][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[20][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[20][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[20][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[20][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[20][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[20][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[20][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[20][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[20][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n112 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[20][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[20][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[20][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[20][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[20][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[21][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[21][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[21][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[21][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[21][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[21][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[21][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[21][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[21][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[21][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[21][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[21][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[21][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[21][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[21][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[21][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[21][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[21][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[21][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[21][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[21][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[21][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[21][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[21][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[21][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[21][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[21][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[21][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[21][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[21][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[21][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[21][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[21][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[21][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[21][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[21][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n111 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[21][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[21][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[21][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[21][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[21][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[22][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[22][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[22][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[22][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[22][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[22][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[22][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[22][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[22][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[22][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[22][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[22][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[22][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[22][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[22][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[22][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[22][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[22][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[22][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[22][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[22][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[22][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[22][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[22][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[22][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[22][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[22][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[22][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[22][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[22][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[22][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[22][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[22][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[22][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[22][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[22][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n110 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[22][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[22][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[22][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[22][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[22][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[23][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[23][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[23][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[23][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[23][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[23][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[23][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[23][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[23][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[23][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[23][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[23][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[23][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[23][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[23][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[23][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[23][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[23][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[23][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[23][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[23][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[23][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[23][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[23][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[23][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[23][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[23][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[23][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[23][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[23][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[23][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[23][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[23][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[23][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[23][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[23][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n109 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[23][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[23][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[23][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[23][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[23][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[24][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[24][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[24][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[24][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[24][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[24][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[24][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[24][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[24][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[24][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[24][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[24][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[24][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[24][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[24][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[24][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[24][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[24][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[24][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[24][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[24][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[24][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[24][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[24][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[24][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[24][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[24][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[24][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[24][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[24][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[24][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[24][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[24][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[24][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[24][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[24][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n108 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[24][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[24][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[24][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[24][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[24][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[25][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[25][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[25][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[25][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[25][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[25][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[25][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[25][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[25][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[25][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[25][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[25][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[25][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[25][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[25][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[25][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[25][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[25][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[25][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[25][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[25][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[25][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[25][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[25][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[25][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[25][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[25][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[25][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[25][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[25][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[25][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[25][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[25][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[25][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[25][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[25][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n107 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[25][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[25][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[25][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[25][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[25][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[26][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[26][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[26][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[26][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[26][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[26][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[26][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[26][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[26][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[26][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[26][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[26][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[26][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[26][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[26][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[26][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[26][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[26][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[26][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[26][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[26][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[26][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[26][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[26][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[26][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[26][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[26][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[26][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[26][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[26][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[26][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[26][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[26][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[26][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[26][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[26][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n106 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[26][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[26][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[26][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[26][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[26][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[27][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[27][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[27][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[27][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[27][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[27][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[27][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[27][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[27][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[27][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[27][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[27][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[27][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[27][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[27][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[27][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[27][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[27][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[27][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[27][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[27][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[27][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[27][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[27][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[27][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[27][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[27][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[27][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[27][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[27][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[27][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[27][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[27][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[27][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[27][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[27][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n105 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[27][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[27][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[27][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[27][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[27][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[28][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[28][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[28][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[28][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[28][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[28][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[28][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[28][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[28][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[28][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[28][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[28][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[28][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[28][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[28][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[28][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[28][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[28][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[28][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[28][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[28][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[28][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[28][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[28][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[28][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[28][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[28][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[28][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[28][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[28][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[28][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[28][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[28][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[28][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[28][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[28][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n104 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[28][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[28][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[28][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[28][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[28][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[29][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[29][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[29][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[29][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[29][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[29][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[29][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[29][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[29][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[29][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[29][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[29][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[29][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[29][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[29][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[29][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[29][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[29][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[29][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[29][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[29][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[29][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[29][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[29][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[29][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[29][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[29][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[29][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[29][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[29][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[29][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[29][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[29][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[29][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[29][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[29][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n103 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[29][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[29][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[29][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[29][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[29][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[30][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[30][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[30][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[30][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[30][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[30][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[30][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[30][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[30][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[30][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[30][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[30][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[30][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[30][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[30][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[30][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[30][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[30][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[30][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[30][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[30][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[30][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[30][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[30][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[30][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[30][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[30][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[30][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[30][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[30][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[30][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[30][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[30][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[30][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[30][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[30][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n102 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[30][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[30][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[30][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[30][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[30][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[31][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[31][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[31][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[31][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[31][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[31][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[31][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[31][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[31][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[31][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[31][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[31][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[31][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[31][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[31][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[31][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[31][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[31][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[31][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[31][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[31][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[31][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[31][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[31][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[31][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[31][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[31][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[31][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[31][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[31][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[31][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[31][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[31][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[31][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[31][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[31][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n101 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[31][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[31][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[31][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[31][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[31][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[32][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[32][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[32][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[32][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[32][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[32][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[32][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[32][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[32][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[32][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[32][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[32][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[32][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[32][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[32][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[32][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[32][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[32][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[32][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[32][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[32][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[32][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[32][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[32][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[32][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[32][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[32][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[32][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[32][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[32][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[32][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[32][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[32][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[32][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[32][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[32][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n100 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[32][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[32][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[32][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[32][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[32][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[33][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[33][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[33][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[33][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[33][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[33][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[33][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[33][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[33][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[33][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[33][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[33][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[33][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[33][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[33][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[33][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[33][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[33][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[33][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[33][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[33][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[33][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[33][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[33][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[33][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[33][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[33][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[33][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[33][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[33][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[33][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[33][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[33][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[33][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[33][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[33][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n99 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[33][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[33][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[33][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[33][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[33][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[34][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[34][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[34][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[34][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[34][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[34][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[34][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[34][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[34][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[34][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[34][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[34][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[34][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[34][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[34][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[34][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[34][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[34][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[34][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[34][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[34][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[34][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[34][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[34][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[34][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[34][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[34][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[34][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[34][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[34][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[34][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[34][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[34][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[34][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[34][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[34][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n98 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[34][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[34][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[34][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[34][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[34][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[35][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[35][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[35][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[35][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[35][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[35][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[35][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[35][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[35][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[35][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[35][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[35][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[35][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[35][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[35][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[35][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[35][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[35][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[35][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[35][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[35][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[35][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[35][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[35][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[35][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[35][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[35][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[35][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[35][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[35][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[35][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[35][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[35][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[35][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[35][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[35][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n97 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[35][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[35][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[35][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[35][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[35][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[36][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[36][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[36][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[36][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[36][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[36][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[36][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[36][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[36][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[36][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[36][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[36][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[36][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[36][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[36][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[36][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[36][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[36][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[36][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[36][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[36][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[36][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[36][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[36][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[36][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[36][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[36][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[36][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[36][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[36][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[36][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[36][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[36][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[36][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[36][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[36][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n96 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[36][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[36][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[36][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[36][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[36][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[37][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[37][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[37][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[37][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[37][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[37][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[37][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[37][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[37][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[37][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[37][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[37][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[37][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[37][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[37][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[37][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[37][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[37][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[37][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[37][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[37][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[37][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[37][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[37][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[37][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[37][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[37][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[37][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[37][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[37][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[37][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[37][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[37][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[37][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[37][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[37][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n95 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[37][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[37][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[37][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[37][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[37][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[38][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[38][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[38][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[38][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[38][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[38][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[38][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[38][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[38][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[38][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[38][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[38][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[38][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[38][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[38][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[38][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[38][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[38][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[38][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[38][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[38][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[38][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[38][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[38][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[38][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[38][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[38][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[38][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[38][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[38][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[38][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[38][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[38][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[38][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[38][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[38][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n94 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[38][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[38][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[38][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[38][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[38][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[39][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[39][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[39][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[39][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[39][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[39][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[39][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[39][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[39][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[39][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[39][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[39][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[39][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[39][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[39][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[39][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[39][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[39][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[39][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[39][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[39][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[39][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[39][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[39][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[39][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[39][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[39][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[39][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[39][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[39][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[39][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[39][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[39][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[39][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[39][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[39][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n93 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[39][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[39][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[39][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[39][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[39][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[40][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[40][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[40][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[40][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[40][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[40][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[40][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[40][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[40][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[40][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[40][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[40][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[40][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[40][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[40][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[40][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[40][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[40][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[40][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[40][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[40][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[40][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[40][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[40][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[40][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[40][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[40][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[40][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[40][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[40][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[40][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[40][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[40][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[40][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[40][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[40][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n92 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[40][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[40][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[40][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[40][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[40][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[41][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[41][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[41][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[41][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[41][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[41][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[41][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[41][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[41][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[41][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[41][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[41][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[41][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[41][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[41][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[41][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[41][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[41][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[41][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[41][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[41][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[41][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[41][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[41][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[41][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[41][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[41][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[41][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[41][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[41][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[41][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[41][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[41][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[41][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[41][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[41][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n91 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[41][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[41][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[41][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[41][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[41][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[42][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[42][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[42][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[42][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[42][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[42][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[42][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[42][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[42][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[42][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[42][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[42][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[42][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[42][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[42][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[42][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[42][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[42][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[42][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[42][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[42][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[42][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[42][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[42][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[42][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[42][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[42][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[42][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[42][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[42][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[42][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[42][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[42][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[42][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[42][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[42][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n90 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[42][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[42][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[42][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[42][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[42][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[43][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[43][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[43][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[43][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[43][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[43][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[43][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[43][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[43][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[43][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[43][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[43][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[43][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[43][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[43][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[43][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[43][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[43][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[43][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[43][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[43][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[43][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[43][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[43][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[43][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[43][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[43][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[43][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[43][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[43][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[43][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[43][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[43][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[43][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[43][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[43][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n89 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[43][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[43][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[43][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[43][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[43][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[44][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[44][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[44][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[44][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[44][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[44][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[44][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[44][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[44][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[44][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[44][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[44][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[44][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[44][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[44][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[44][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[44][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[44][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[44][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[44][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[44][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[44][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[44][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[44][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[44][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[44][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[44][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[44][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[44][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[44][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[44][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[44][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[44][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[44][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[44][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[44][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n88 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[44][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[44][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[44][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[44][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[44][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[45][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[45][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[45][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[45][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[45][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[45][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[45][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[45][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[45][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[45][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[45][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[45][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[45][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[45][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[45][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[45][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[45][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[45][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[45][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[45][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[45][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[45][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[45][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[45][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[45][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[45][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[45][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[45][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[45][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[45][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[45][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[45][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[45][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[45][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[45][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[45][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n87 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[45][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[45][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[45][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[45][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[45][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[46][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[46][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[46][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[46][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[46][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[46][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[46][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[46][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[46][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[46][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[46][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[46][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[46][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[46][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[46][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[46][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[46][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[46][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[46][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[46][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[46][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[46][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[46][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[46][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[46][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[46][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[46][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[46][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[46][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[46][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[46][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[46][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[46][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[46][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[46][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[46][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n86 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[46][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[46][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[46][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[46][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[46][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[47][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[47][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[47][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[47][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[47][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[47][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[47][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[47][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[47][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[47][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[47][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[47][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[47][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[47][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[47][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[47][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[47][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[47][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[47][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[47][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[47][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[47][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[47][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[47][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[47][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[47][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[47][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[47][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[47][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[47][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[47][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[47][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[47][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[47][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[47][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[47][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n85 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[47][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[47][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[47][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[47][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[47][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[48][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[48][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[48][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[48][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[48][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[48][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[48][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[48][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[48][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[48][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[48][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[48][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[48][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[48][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[48][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[48][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[48][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[48][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[48][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[48][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[48][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[48][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[48][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[48][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[48][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[48][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[48][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[48][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[48][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[48][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[48][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[48][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[48][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[48][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[48][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[48][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n84 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[48][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[48][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[48][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[48][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[48][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[49][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[49][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[49][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[49][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[49][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[49][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[49][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[49][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[49][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[49][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[49][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[49][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[49][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[49][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[49][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[49][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[49][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[49][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[49][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[49][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[49][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[49][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[49][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[49][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[49][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[49][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[49][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[49][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[49][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[49][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[49][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[49][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[49][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[49][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[49][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[49][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n83 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[49][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[49][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[49][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[49][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[49][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[50][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[50][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[50][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[50][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[50][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[50][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[50][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[50][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[50][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[50][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[50][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[50][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[50][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[50][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[50][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[50][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[50][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[50][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[50][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[50][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[50][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[50][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[50][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[50][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[50][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[50][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[50][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[50][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[50][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[50][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[50][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[50][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[50][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[50][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[50][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[50][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n82 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[50][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[50][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[50][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[50][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[50][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[51][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[51][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[51][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[51][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[51][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[51][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[51][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[51][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[51][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[51][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[51][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[51][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[51][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[51][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[51][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[51][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[51][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[51][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[51][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[51][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[51][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[51][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[51][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[51][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[51][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[51][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[51][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[51][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[51][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[51][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[51][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[51][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[51][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[51][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[51][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[51][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n81 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[51][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[51][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[51][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[51][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[51][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[52][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[52][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[52][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[52][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[52][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[52][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[52][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[52][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[52][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[52][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[52][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[52][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[52][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[52][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[52][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[52][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[52][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[52][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[52][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[52][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[52][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[52][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[52][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[52][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[52][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[52][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[52][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[52][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[52][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[52][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[52][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[52][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[52][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[52][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[52][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[52][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n80 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[52][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[52][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[52][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[52][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[52][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[53][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[53][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[53][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[53][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[53][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[53][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[53][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[53][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[53][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[53][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[53][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[53][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[53][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[53][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[53][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[53][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[53][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[53][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[53][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[53][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[53][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[53][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[53][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[53][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[53][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[53][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[53][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[53][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[53][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[53][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[53][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[53][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[53][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[53][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[53][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[53][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n79 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[53][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[53][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[53][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[53][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[53][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[54][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[54][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[54][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[54][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[54][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[54][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[54][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[54][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[54][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[54][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[54][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[54][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[54][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[54][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[54][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[54][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[54][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[54][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[54][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[54][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[54][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[54][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[54][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[54][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[54][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[54][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[54][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[54][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[54][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[54][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[54][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[54][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[54][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[54][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[54][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[54][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n78 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[54][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[54][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[54][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[54][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[54][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[55][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[55][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[55][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[55][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[55][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[55][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[55][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[55][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[55][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[55][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[55][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[55][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[55][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[55][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[55][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[55][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[55][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[55][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[55][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[55][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[55][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[55][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[55][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[55][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[55][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[55][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[55][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[55][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[55][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[55][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[55][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[55][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[55][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[55][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[55][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[55][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n77 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[55][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[55][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[55][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[55][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[55][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[56][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[56][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[56][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[56][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[56][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[56][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[56][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[56][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[56][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[56][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[56][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[56][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[56][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[56][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[56][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[56][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[56][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[56][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[56][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[56][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[56][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[56][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[56][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[56][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[56][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[56][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[56][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[56][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[56][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[56][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[56][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[56][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[56][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[56][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[56][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[56][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n76 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[56][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[56][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[56][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[56][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[56][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[57][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[57][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[57][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[57][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[57][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[57][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[57][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[57][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[57][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[57][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[57][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[57][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[57][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[57][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[57][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[57][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[57][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[57][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[57][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[57][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[57][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[57][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[57][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[57][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[57][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[57][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[57][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[57][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[57][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[57][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[57][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[57][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[57][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[57][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[57][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[57][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n75 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[57][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[57][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[57][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[57][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[57][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[58][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[58][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[58][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[58][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[58][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[58][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[58][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[58][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[58][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[58][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[58][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[58][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[58][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[58][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[58][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[58][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[58][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[58][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[58][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[58][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[58][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[58][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[58][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[58][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[58][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[58][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[58][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[58][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[58][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[58][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[58][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[58][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[58][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[58][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[58][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[58][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n74 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[58][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[58][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[58][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[58][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[58][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[59][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[59][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[59][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[59][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[59][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[59][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[59][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[59][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[59][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[59][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[59][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[59][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[59][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[59][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[59][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[59][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[59][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[59][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[59][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[59][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[59][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[59][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[59][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[59][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[59][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[59][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[59][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[59][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[59][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[59][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[59][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[59][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[59][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[59][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[59][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[59][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n73 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[59][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[59][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[59][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[59][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[59][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[60][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[60][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[60][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[60][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[60][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[60][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[60][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[60][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[60][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[60][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[60][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[60][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[60][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[60][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[60][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[60][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[60][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[60][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[60][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[60][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[60][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[60][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[60][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[60][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[60][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[60][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[60][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[60][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[60][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[60][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[60][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[60][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[60][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[60][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[60][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[60][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n72 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[60][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[60][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[60][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[60][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[60][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[61][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[61][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[61][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[61][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[61][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[61][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[61][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[61][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[61][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[61][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[61][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[61][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[61][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[61][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[61][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[61][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[61][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[61][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[61][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[61][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[61][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[61][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[61][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[61][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[61][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[61][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[61][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[61][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[61][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[61][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[61][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[61][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[61][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[61][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[61][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[61][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n71 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[61][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[61][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[61][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[61][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[61][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[62][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[62][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[62][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[62][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[62][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[62][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[62][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[62][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[62][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[62][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[62][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[62][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[62][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[62][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[62][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[62][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[62][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[62][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[62][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[62][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[62][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[62][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[62][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[62][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[62][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[62][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[62][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[62][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[62][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[62][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[62][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[62][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[62][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[62][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[62][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[62][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n70 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[62][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[62][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[62][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[62][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[62][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[63][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[63][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[63][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[63][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[63][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[63][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[63][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[63][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[63][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[63][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[63][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[63][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[63][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[63][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[63][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[63][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[63][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[63][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[63][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[63][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[63][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[63][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[63][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[63][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[63][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[63][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[63][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[63][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[63][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[63][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[63][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[63][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[63][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[63][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[63][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[63][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n69 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[63][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[63][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[63][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[63][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[63][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[64][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[64][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[64][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[64][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[64][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[64][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[64][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[64][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[64][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[64][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[64][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[64][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[64][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[64][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[64][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[64][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[64][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[64][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[64][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[64][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[64][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[64][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[64][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[64][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[64][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[64][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[64][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[64][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[64][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[64][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[64][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[64][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[64][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[64][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[64][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[64][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n68 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[64][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[64][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[64][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[64][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[64][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[65][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[65][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[65][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[65][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[65][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[65][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[65][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[65][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[65][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[65][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[65][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[65][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[65][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[65][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[65][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[65][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[65][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[65][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[65][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[65][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[65][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[65][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[65][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[65][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[65][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[65][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[65][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[65][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[65][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[65][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[65][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[65][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[65][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[65][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[65][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[65][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n67 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[65][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[65][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[65][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[65][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[65][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[66][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[66][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[66][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[66][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[66][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[66][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[66][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[66][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[66][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[66][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[66][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[66][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[66][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[66][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[66][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[66][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[66][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[66][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[66][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[66][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[66][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[66][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[66][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[66][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[66][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[66][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[66][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[66][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[66][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[66][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[66][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[66][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[66][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[66][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[66][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[66][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n66 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[66][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[66][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[66][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[66][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[66][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[67][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[67][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[67][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[67][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[67][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[67][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[67][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[67][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[67][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[67][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[67][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[67][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[67][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[67][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[67][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[67][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[67][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[67][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[67][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[67][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[67][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[67][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[67][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[67][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[67][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[67][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[67][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[67][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[67][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[67][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[67][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[67][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[67][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[67][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[67][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[67][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n65 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[67][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[67][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[67][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[67][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[67][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[68][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[68][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[68][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[68][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[68][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[68][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[68][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[68][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[68][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[68][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[68][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[68][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[68][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[68][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[68][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[68][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[68][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[68][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[68][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[68][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[68][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[68][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[68][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[68][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[68][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[68][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[68][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[68][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[68][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[68][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[68][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[68][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[68][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[68][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[68][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[68][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n64 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[68][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[68][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[68][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[68][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[68][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[69][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[69][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[69][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[69][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[69][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[69][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[69][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[69][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[69][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[69][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[69][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[69][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[69][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[69][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[69][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[69][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[69][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[69][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[69][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[69][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[69][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[69][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[69][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[69][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[69][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[69][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[69][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[69][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[69][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[69][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[69][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[69][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[69][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[69][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[69][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[69][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n63 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[69][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[69][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[69][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[69][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[69][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[70][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[70][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[70][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[70][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[70][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[70][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[70][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[70][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[70][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[70][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[70][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[70][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[70][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[70][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[70][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[70][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[70][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[70][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[70][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[70][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[70][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[70][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[70][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[70][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[70][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[70][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[70][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[70][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[70][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[70][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[70][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[70][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[70][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[70][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[70][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[70][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n62 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[70][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[70][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[70][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[70][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[70][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[71][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[71][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[71][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[71][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[71][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[71][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[71][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[71][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[71][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[71][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[71][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[71][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[71][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[71][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[71][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[71][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[71][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[71][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[71][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[71][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[71][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[71][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[71][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[71][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[71][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[71][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[71][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[71][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[71][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[71][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[71][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[71][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[71][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[71][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[71][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[71][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n61 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[71][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[71][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[71][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[71][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[71][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[72][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[72][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[72][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[72][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[72][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[72][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[72][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[72][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[72][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[72][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[72][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[72][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[72][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[72][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[72][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[72][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[72][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[72][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[72][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[72][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[72][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[72][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[72][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[72][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[72][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[72][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[72][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[72][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[72][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[72][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[72][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[72][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[72][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[72][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[72][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[72][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n60 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[72][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[72][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[72][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[72][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[72][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[73][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[73][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[73][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[73][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[73][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[73][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[73][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[73][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[73][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[73][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[73][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[73][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[73][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[73][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[73][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[73][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[73][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[73][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[73][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[73][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[73][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[73][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[73][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[73][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[73][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[73][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[73][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[73][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[73][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[73][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[73][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[73][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[73][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[73][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[73][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[73][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n59 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[73][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[73][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[73][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[73][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[73][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[74][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[74][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[74][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[74][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[74][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[74][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[74][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[74][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[74][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[74][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[74][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[74][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[74][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[74][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[74][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[74][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[74][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[74][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[74][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[74][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[74][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[74][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[74][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[74][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[74][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[74][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[74][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[74][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[74][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[74][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[74][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[74][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[74][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[74][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[74][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[74][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n58 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[74][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[74][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[74][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[74][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[74][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[75][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[75][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[75][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[75][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[75][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[75][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[75][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[75][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[75][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[75][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[75][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[75][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[75][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[75][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[75][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[75][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[75][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[75][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[75][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[75][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[75][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[75][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[75][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[75][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[75][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[75][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[75][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[75][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[75][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[75][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[75][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[75][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[75][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[75][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[75][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[75][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n57 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[75][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[75][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[75][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[75][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[75][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[76][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[76][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[76][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[76][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[76][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[76][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[76][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[76][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[76][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[76][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[76][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[76][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[76][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[76][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[76][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[76][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[76][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[76][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[76][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[76][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[76][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[76][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[76][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[76][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[76][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[76][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[76][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[76][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[76][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[76][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[76][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[76][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[76][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[76][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[76][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[76][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n56 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[76][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[76][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[76][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[76][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[76][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[77][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[77][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[77][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[77][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[77][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[77][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[77][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[77][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[77][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[77][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[77][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[77][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[77][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[77][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[77][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[77][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[77][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[77][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[77][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[77][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[77][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[77][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[77][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[77][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[77][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[77][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[77][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[77][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[77][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[77][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[77][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[77][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[77][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[77][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[77][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[77][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n55 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[77][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[77][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[77][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[77][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[77][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[78][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[78][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[78][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[78][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[78][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[78][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[78][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[78][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[78][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[78][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[78][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[78][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[78][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[78][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[78][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[78][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[78][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[78][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[78][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[78][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[78][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[78][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[78][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[78][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[78][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[78][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[78][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[78][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[78][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[78][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[78][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[78][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[78][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[78][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[78][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[78][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n54 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[78][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[78][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[78][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[78][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[78][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[79][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[79][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[79][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[79][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[79][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[79][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[79][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[79][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[79][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[79][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[79][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[79][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[79][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[79][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[79][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[79][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[79][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[79][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[79][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[79][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[79][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[79][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[79][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[79][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[79][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[79][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[79][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[79][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[79][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[79][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[79][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[79][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[79][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[79][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[79][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[79][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n53 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[79][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[79][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[79][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[79][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[79][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[80][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[80][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[80][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[80][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[80][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[80][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[80][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[80][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[80][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[80][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[80][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[80][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[80][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[80][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[80][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[80][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[80][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[80][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[80][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[80][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[80][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[80][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[80][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[80][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[80][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[80][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[80][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[80][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[80][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[80][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[80][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[80][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[80][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[80][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[80][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[80][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n52 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[80][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[80][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[80][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[80][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[80][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[81][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[81][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[81][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[81][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[81][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[81][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[81][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[81][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[81][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[81][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[81][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[81][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[81][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[81][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[81][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[81][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[81][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[81][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[81][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[81][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[81][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[81][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[81][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[81][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[81][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[81][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[81][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[81][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[81][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[81][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[81][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[81][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[81][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[81][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[81][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[81][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n51 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[81][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[81][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[81][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[81][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[81][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[82][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[82][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[82][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[82][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[82][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[82][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[82][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[82][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[82][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[82][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[82][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[82][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[82][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[82][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[82][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[82][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[82][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[82][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[82][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[82][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[82][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[82][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[82][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[82][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[82][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[82][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[82][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[82][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[82][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[82][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[82][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[82][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[82][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[82][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[82][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[82][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n50 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[82][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[82][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[82][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[82][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[82][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[83][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[83][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[83][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[83][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[83][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[83][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[83][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[83][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[83][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[83][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[83][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[83][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[83][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[83][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[83][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[83][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[83][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[83][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[83][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[83][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[83][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[83][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[83][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[83][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[83][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[83][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[83][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[83][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[83][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[83][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[83][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[83][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[83][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[83][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[83][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[83][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n49 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[83][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[83][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[83][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[83][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[83][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[84][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[84][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[84][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[84][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[84][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[84][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[84][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[84][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[84][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[84][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[84][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[84][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[84][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[84][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[84][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[84][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[84][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[84][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[84][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[84][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[84][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[84][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[84][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[84][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[84][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[84][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[84][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[84][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[84][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[84][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[84][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[84][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[84][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[84][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[84][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[84][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n48 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[84][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[84][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[84][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[84][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[84][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[85][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[85][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[85][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[85][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[85][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[85][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[85][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[85][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[85][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[85][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[85][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[85][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[85][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[85][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[85][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[85][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[85][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[85][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[85][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[85][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[85][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[85][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[85][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[85][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[85][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[85][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[85][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[85][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[85][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[85][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[85][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[85][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[85][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[85][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[85][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[85][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n47 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[85][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[85][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[85][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[85][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[85][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[86][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[86][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[86][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[86][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[86][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[86][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[86][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[86][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[86][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[86][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[86][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[86][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[86][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[86][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[86][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[86][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[86][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[86][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[86][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[86][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[86][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[86][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[86][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[86][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[86][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[86][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[86][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[86][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[86][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[86][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[86][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[86][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[86][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[86][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[86][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[86][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n46 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[86][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[86][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[86][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[86][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[86][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[87][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[87][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[87][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[87][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[87][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[87][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[87][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[87][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[87][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[87][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[87][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[87][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[87][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[87][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[87][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[87][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[87][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[87][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[87][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[87][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[87][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[87][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[87][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[87][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[87][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[87][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[87][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[87][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[87][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[87][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[87][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[87][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[87][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[87][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[87][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[87][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n45 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[87][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[87][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[87][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[87][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[87][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[88][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[88][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[88][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[88][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[88][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[88][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[88][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[88][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[88][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[88][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[88][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[88][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[88][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[88][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[88][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[88][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[88][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[88][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[88][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[88][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[88][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[88][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[88][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[88][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[88][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[88][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[88][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[88][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[88][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[88][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[88][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[88][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[88][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[88][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[88][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[88][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n44 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[88][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[88][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[88][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[88][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[88][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[89][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[89][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[89][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[89][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[89][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[89][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[89][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[89][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[89][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[89][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[89][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[89][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[89][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[89][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[89][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[89][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[89][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[89][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[89][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[89][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[89][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[89][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[89][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[89][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[89][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[89][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[89][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[89][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[89][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[89][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[89][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[89][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[89][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[89][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[89][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[89][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n43 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[89][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[89][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[89][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[89][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[89][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[90][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[90][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[90][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[90][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[90][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[90][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[90][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[90][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[90][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[90][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[90][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[90][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[90][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[90][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[90][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[90][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[90][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[90][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[90][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[90][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[90][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[90][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[90][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[90][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[90][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[90][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[90][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[90][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[90][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[90][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[90][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[90][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[90][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[90][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[90][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[90][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n42 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[90][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[90][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[90][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[90][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[90][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[91][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[91][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[91][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[91][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[91][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[91][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[91][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[91][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[91][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[91][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[91][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[91][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[91][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[91][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[91][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[91][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[91][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[91][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[91][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[91][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[91][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[91][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[91][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[91][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[91][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[91][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[91][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[91][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[91][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[91][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[91][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[91][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[91][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[91][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[91][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[91][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n41 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[91][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[91][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[91][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[91][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[91][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[92][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[92][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[92][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[92][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[92][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[92][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[92][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[92][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[92][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[92][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[92][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[92][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[92][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[92][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[92][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[92][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[92][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[92][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[92][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[92][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[92][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[92][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[92][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[92][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[92][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[92][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[92][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[92][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[92][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[92][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[92][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[92][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[92][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[92][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[92][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[92][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n40 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[92][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[92][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[92][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[92][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[92][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[93][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[93][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[93][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[93][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[93][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[93][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[93][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[93][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[93][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[93][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[93][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[93][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[93][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[93][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[93][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[93][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[93][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[93][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[93][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[93][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[93][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[93][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[93][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[93][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[93][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[93][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[93][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[93][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[93][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[93][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[93][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[93][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[93][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[93][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[93][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[93][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n39 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[93][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[93][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[93][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[93][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[93][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[94][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[94][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[94][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[94][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[94][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[94][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[94][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[94][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[94][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[94][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[94][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[94][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[94][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[94][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[94][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[94][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[94][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[94][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[94][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[94][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[94][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[94][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[94][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[94][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[94][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[94][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[94][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[94][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[94][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[94][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[94][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[94][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[94][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[94][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[94][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[94][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n38 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[94][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[94][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[94][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[94][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[94][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[95][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[95][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[95][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[95][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[95][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[95][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[95][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[95][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[95][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[95][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[95][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[95][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[95][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[95][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[95][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[95][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[95][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[95][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[95][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[95][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[95][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[95][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[95][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[95][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[95][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[95][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[95][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[95][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[95][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[95][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[95][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[95][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[95][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[95][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[95][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[95][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n37 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[95][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[95][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[95][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[95][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[95][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[96][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[96][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[96][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[96][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[96][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[96][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[96][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[96][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[96][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[96][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[96][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[96][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[96][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[96][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[96][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[96][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[96][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[96][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[96][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[96][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[96][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[96][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[96][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[96][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[96][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[96][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[96][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[96][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[96][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[96][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[96][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[96][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[96][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[96][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[96][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[96][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n36 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[96][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[96][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[96][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[96][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[96][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[97][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[97][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[97][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[97][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[97][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[97][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[97][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[97][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[97][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[97][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[97][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[97][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[97][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[97][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[97][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[97][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[97][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[97][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[97][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[97][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[97][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[97][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[97][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[97][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[97][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[97][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[97][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[97][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[97][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[97][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[97][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[97][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[97][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[97][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[97][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[97][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n35 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[97][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[97][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[97][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[97][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[97][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[98][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[98][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[98][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[98][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[98][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[98][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[98][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[98][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[98][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[98][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[98][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[98][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[98][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[98][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[98][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[98][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[98][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[98][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[98][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[98][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[98][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[98][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[98][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[98][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[98][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[98][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[98][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[98][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[98][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[98][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[98][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[98][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[98][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[98][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[98][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[98][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n34 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[98][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[98][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[98][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[98][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[98][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[99][0]~FF  (.D(\data_to_rx_packet_reg[0] ), .CE(\i16/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[99][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[99][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[99][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[99][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[99][1]~FF  (.D(\data_to_rx_packet_reg[1] ), .CE(\i16/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[99][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[99][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[99][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[99][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[99][2]~FF  (.D(\data_to_rx_packet_reg[2] ), .CE(\i16/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[99][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[99][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[99][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[99][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[99][3]~FF  (.D(\data_to_rx_packet_reg[3] ), .CE(\i16/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[99][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[99][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[99][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[99][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[99][4]~FF  (.D(\data_to_rx_packet_reg[4] ), .CE(\i16/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[99][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[99][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[99][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[99][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[99][5]~FF  (.D(\data_to_rx_packet_reg[5] ), .CE(\i16/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[99][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[99][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[99][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[99][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[99][6]~FF  (.D(\data_to_rx_packet_reg[6] ), .CE(\i16/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[99][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[99][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[99][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[99][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[99][7]~FF  (.D(\data_to_rx_packet_reg[7] ), .CE(\i16/n33 ), 
           .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[99][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[99][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[99][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[99][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[99][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[100][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[100][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[100][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[100][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[100][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[100][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[100][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[100][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[100][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[100][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[100][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[100][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[100][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[100][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[100][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[100][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[100][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[100][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[100][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[100][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[100][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[100][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[100][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[100][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[100][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[100][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[100][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[100][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[100][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[100][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[100][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[100][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[100][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[100][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[100][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[100][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n32 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[100][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[100][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[100][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[100][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[100][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[101][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[101][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[101][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[101][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[101][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[101][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[101][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[101][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[101][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[101][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[101][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[101][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[101][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[101][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[101][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[101][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[101][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[101][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[101][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[101][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[101][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[101][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[101][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[101][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[101][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[101][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[101][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[101][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[101][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[101][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[101][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[101][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[101][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[101][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[101][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[101][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n31 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[101][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[101][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[101][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[101][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[101][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[102][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[102][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[102][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[102][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[102][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[102][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[102][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[102][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[102][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[102][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[102][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[102][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[102][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[102][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[102][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[102][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[102][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[102][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[102][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[102][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[102][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[102][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[102][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[102][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[102][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[102][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[102][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[102][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[102][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[102][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[102][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[102][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[102][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[102][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[102][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[102][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n30 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[102][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[102][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[102][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[102][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[102][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[103][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[103][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[103][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[103][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[103][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[103][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[103][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[103][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[103][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[103][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[103][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[103][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[103][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[103][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[103][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[103][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[103][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[103][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[103][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[103][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[103][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[103][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[103][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[103][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[103][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[103][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[103][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[103][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[103][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[103][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[103][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[103][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[103][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[103][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[103][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[103][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n29 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[103][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[103][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[103][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[103][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[103][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[104][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[104][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[104][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[104][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[104][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[104][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[104][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[104][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[104][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[104][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[104][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[104][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[104][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[104][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[104][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[104][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[104][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[104][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[104][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[104][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[104][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[104][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[104][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[104][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[104][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[104][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[104][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[104][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[104][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[104][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[104][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[104][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[104][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[104][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[104][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[104][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n28 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[104][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[104][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[104][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[104][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[104][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[105][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[105][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[105][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[105][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[105][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[105][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[105][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[105][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[105][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[105][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[105][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[105][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[105][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[105][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[105][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[105][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[105][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[105][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[105][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[105][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[105][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[105][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[105][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[105][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[105][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[105][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[105][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[105][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[105][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[105][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[105][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[105][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[105][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[105][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[105][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[105][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n27 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[105][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[105][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[105][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[105][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[105][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[106][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[106][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[106][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[106][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[106][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[106][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[106][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[106][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[106][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[106][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[106][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[106][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[106][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[106][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[106][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[106][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[106][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[106][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[106][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[106][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[106][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[106][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[106][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[106][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[106][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[106][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[106][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[106][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[106][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[106][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[106][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[106][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[106][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[106][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[106][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[106][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n26 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[106][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[106][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[106][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[106][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[106][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[107][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[107][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[107][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[107][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[107][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[107][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[107][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[107][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[107][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[107][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[107][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[107][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[107][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[107][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[107][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[107][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[107][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[107][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[107][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[107][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[107][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[107][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[107][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[107][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[107][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[107][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[107][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[107][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[107][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[107][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[107][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[107][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[107][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[107][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[107][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[107][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n25 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[107][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[107][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[107][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[107][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[107][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[108][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[108][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[108][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[108][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[108][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[108][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[108][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[108][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[108][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[108][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[108][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[108][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[108][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[108][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[108][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[108][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[108][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[108][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[108][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[108][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[108][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[108][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[108][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[108][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[108][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[108][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[108][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[108][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[108][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[108][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[108][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[108][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[108][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[108][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[108][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[108][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n24 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[108][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[108][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[108][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[108][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[108][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[109][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[109][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[109][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[109][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[109][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[109][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[109][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[109][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[109][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[109][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[109][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[109][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[109][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[109][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[109][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[109][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[109][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[109][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[109][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[109][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[109][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[109][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[109][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[109][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[109][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[109][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[109][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[109][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[109][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[109][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[109][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[109][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[109][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[109][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[109][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[109][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n23 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[109][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[109][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[109][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[109][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[109][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[110][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[110][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[110][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[110][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[110][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[110][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[110][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[110][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[110][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[110][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[110][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[110][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[110][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[110][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[110][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[110][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[110][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[110][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[110][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[110][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[110][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[110][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[110][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[110][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[110][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[110][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[110][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[110][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[110][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[110][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[110][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[110][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[110][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[110][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[110][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[110][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n22 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[110][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[110][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[110][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[110][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[110][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[111][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[111][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[111][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[111][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[111][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[111][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[111][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[111][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[111][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[111][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[111][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[111][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[111][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[111][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[111][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[111][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[111][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[111][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[111][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[111][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[111][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[111][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[111][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[111][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[111][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[111][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[111][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[111][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[111][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[111][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[111][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[111][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[111][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[111][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[111][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[111][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n21 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[111][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[111][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[111][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[111][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[111][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[112][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[112][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[112][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[112][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[112][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[112][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[112][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[112][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[112][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[112][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[112][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[112][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[112][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[112][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[112][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[112][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[112][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[112][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[112][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[112][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[112][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[112][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[112][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[112][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[112][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[112][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[112][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[112][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[112][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[112][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[112][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[112][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[112][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[112][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[112][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[112][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n20 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[112][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[112][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[112][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[112][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[112][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[113][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[113][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[113][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[113][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[113][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[113][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[113][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[113][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[113][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[113][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[113][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[113][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[113][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[113][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[113][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[113][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[113][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[113][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[113][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[113][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[113][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[113][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[113][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[113][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[113][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[113][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[113][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[113][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[113][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[113][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[113][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[113][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[113][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[113][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[113][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[113][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n19 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[113][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[113][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[113][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[113][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[113][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[114][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[114][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[114][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[114][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[114][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[114][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[114][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[114][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[114][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[114][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[114][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[114][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[114][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[114][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[114][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[114][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[114][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[114][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[114][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[114][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[114][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[114][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[114][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[114][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[114][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[114][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[114][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[114][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[114][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[114][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[114][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[114][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[114][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[114][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[114][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[114][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n18 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[114][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[114][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[114][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[114][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[114][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[115][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[115][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[115][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[115][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[115][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[115][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[115][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[115][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[115][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[115][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[115][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[115][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[115][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[115][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[115][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[115][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[115][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[115][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[115][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[115][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[115][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[115][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[115][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[115][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[115][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[115][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[115][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[115][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[115][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[115][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[115][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[115][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[115][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[115][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[115][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[115][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n17 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[115][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[115][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[115][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[115][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[115][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[116][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[116][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[116][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[116][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[116][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[116][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[116][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[116][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[116][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[116][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[116][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[116][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[116][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[116][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[116][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[116][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[116][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[116][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[116][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[116][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[116][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[116][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[116][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[116][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[116][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[116][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[116][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[116][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[116][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[116][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[116][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[116][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[116][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[116][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[116][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[116][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n16 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[116][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[116][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[116][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[116][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[116][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[117][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[117][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[117][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[117][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[117][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[117][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[117][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[117][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[117][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[117][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[117][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[117][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[117][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[117][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[117][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[117][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[117][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[117][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[117][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[117][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[117][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[117][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[117][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[117][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[117][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[117][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[117][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[117][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[117][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[117][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[117][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[117][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[117][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[117][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[117][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[117][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n15 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[117][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[117][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[117][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[117][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[117][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[118][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[118][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[118][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[118][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[118][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[118][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[118][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[118][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[118][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[118][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[118][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[118][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[118][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[118][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[118][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[118][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[118][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[118][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[118][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[118][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[118][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[118][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[118][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[118][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[118][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[118][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[118][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[118][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[118][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[118][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[118][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[118][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[118][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[118][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[118][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[118][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n14 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[118][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[118][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[118][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[118][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[118][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[119][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[119][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[119][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[119][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[119][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[119][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[119][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[119][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[119][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[119][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[119][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[119][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[119][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[119][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[119][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[119][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[119][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[119][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[119][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[119][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[119][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[119][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[119][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[119][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[119][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[119][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[119][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[119][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[119][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[119][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[119][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[119][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[119][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[119][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[119][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[119][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n13 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[119][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[119][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[119][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[119][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[119][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[120][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[120][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[120][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[120][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[120][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[120][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[120][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[120][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[120][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[120][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[120][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[120][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[120][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[120][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[120][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[120][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[120][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[120][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[120][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[120][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[120][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[120][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[120][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[120][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[120][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[120][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[120][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[120][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[120][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[120][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[120][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[120][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[120][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[120][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[120][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[120][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n12 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[120][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[120][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[120][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[120][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[120][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[121][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[121][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[121][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[121][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[121][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[121][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[121][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[121][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[121][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[121][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[121][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[121][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[121][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[121][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[121][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[121][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[121][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[121][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[121][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[121][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[121][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[121][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[121][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[121][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[121][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[121][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[121][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[121][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[121][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[121][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[121][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[121][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[121][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[121][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[121][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[121][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n11 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[121][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[121][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[121][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[121][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[121][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[122][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[122][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[122][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[122][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[122][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[122][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[122][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[122][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[122][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[122][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[122][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[122][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[122][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[122][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[122][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[122][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[122][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[122][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[122][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[122][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[122][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[122][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[122][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[122][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[122][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[122][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[122][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[122][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[122][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[122][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[122][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[122][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[122][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[122][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[122][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[122][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n10 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[122][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[122][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[122][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[122][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[122][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[123][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[123][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[123][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[123][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[123][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[123][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[123][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[123][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[123][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[123][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[123][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[123][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[123][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[123][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[123][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[123][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[123][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[123][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[123][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[123][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[123][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[123][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[123][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[123][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[123][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[123][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[123][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[123][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[123][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[123][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[123][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[123][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[123][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[123][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[123][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[123][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n9 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[123][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[123][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[123][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[123][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[123][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[124][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[124][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[124][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[124][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[124][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[124][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[124][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[124][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[124][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[124][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[124][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[124][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[124][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[124][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[124][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[124][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[124][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[124][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[124][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[124][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[124][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[124][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[124][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[124][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[124][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[124][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[124][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[124][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[124][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[124][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[124][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[124][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[124][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[124][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[124][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[124][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n8 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[124][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[124][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[124][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[124][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[124][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[125][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[125][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[125][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[125][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[125][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[125][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[125][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[125][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[125][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[125][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[125][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[125][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[125][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[125][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[125][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[125][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[125][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[125][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[125][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[125][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[125][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[125][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[125][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[125][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[125][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[125][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[125][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[125][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[125][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[125][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[125][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[125][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[125][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[125][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[125][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[125][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n7 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[125][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[125][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[125][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[125][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[125][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[126][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[126][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[126][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[126][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[126][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[126][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[126][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[126][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[126][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[126][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[126][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[126][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[126][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[126][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[126][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[126][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[126][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[126][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[126][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[126][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[126][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[126][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[126][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[126][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[126][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[126][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[126][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[126][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[126][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[126][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[126][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[126][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[126][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[126][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[126][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[126][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n6 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[126][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[126][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[126][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[126][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[126][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[127][0]~FF  (.D(\data_to_rx_packet_reg[0] ), 
           .CE(\i16/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[127][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[127][0]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][0]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][0]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][0]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][0]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[127][0]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[127][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[127][1]~FF  (.D(\data_to_rx_packet_reg[1] ), 
           .CE(\i16/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[127][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[127][1]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][1]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][1]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][1]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][1]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[127][1]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[127][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[127][2]~FF  (.D(\data_to_rx_packet_reg[2] ), 
           .CE(\i16/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[127][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[127][2]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][2]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][2]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][2]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][2]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[127][2]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[127][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[127][3]~FF  (.D(\data_to_rx_packet_reg[3] ), 
           .CE(\i16/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[127][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[127][3]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][3]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][3]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][3]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][3]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[127][3]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[127][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[127][4]~FF  (.D(\data_to_rx_packet_reg[4] ), 
           .CE(\i16/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[127][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[127][4]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][4]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][4]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][4]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][4]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[127][4]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[127][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[127][5]~FF  (.D(\data_to_rx_packet_reg[5] ), 
           .CE(\i16/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[127][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[127][5]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][5]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][5]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][5]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][5]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[127][5]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[127][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[127][6]~FF  (.D(\data_to_rx_packet_reg[6] ), 
           .CE(\i16/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[127][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[127][6]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][6]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][6]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][6]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][6]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[127][6]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[127][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i16/rx_fifo/buff[127][7]~FF  (.D(\data_to_rx_packet_reg[7] ), 
           .CE(\i16/n5 ), .CLK(\pll_clk~O ), .SR(1'b0), .Q(\i16/rx_fifo/buff[127][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(16)
    defparam \i16/rx_fifo/buff[127][7]~FF .CLK_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][7]~FF .CE_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][7]~FF .SR_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][7]~FF .D_POLARITY = 1'b1;
    defparam \i16/rx_fifo/buff[127][7]~FF .SR_SYNC = 1'b1;
    defparam \i16/rx_fifo/buff[127][7]~FF .SR_VALUE = 1'b0;
    defparam \i16/rx_fifo/buff[127][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \tx_dac_fsm_inst/i119  (.I0(n3564), .I1(n115), .I2(n3562), 
            .O(n115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/i119 .LUTMASK = 16'hacac;
    EFX_LUT4 \tx_dac_fsm_inst/dlatchrs_164/i1  (.I0(n3565), .I1(n116), .I2(n3562), 
            .O(n116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/dlatchrs_164/i1 .LUTMASK = 16'hacac;
    EFX_LUT4 \tx_dac_fsm_inst/dlatchrs_162/i2  (.I0(n3583), .I1(n133), .I2(n3557), 
            .O(n133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/dlatchrs_162/i2 .LUTMASK = 16'hacac;
    EFX_LUT4 \tx_dac_fsm_inst/dlatchrs_162/i3  (.I0(n3584), .I1(n134), .I2(n3557), 
            .O(n134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/dlatchrs_162/i3 .LUTMASK = 16'hacac;
    EFX_LUT4 \tx_dac_fsm_inst/dlatchrs_162/i4  (.I0(n3585), .I1(n135), .I2(n3557), 
            .O(n135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/dlatchrs_162/i4 .LUTMASK = 16'hacac;
    EFX_LUT4 \tx_dac_fsm_inst/dlatchrs_164/i2  (.I0(n3586), .I1(n136), .I2(n3562), 
            .O(n136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/dlatchrs_164/i2 .LUTMASK = 16'hacac;
    EFX_LUT4 LUT__7662 (.I0(\spi_slave_inst/bitcnt[4] ), .I1(\spi_slave_inst/bitcnt[3] ), 
            .O(n4235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7662.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7663 (.I0(n4235), .I1(rw_out), .I2(\spi_slave_inst/d_o[7] ), 
            .O(MISO)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__7663.LUTMASK = 16'h4040;
    EFX_ADD \led_inst/add_23/i2  (.I0(\led_inst/counter[1] ), .I1(\led_inst/counter[0] ), 
            .CI(1'b0), .O(n19), .CO(n20)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i2 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_129/i2  (.I0(\tx_dac_fsm_inst/zctr[1] ), 
            .I1(\tx_dac_fsm_inst/zctr[0] ), .CI(1'b0), .O(n118), .CO(n119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(197)
    defparam \tx_dac_fsm_inst/add_129/i2 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_129/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_136/i2  (.I0(\tx_dac_fsm_inst/dctr[1] ), 
            .I1(\tx_dac_fsm_inst/dctr[0] ), .CI(1'b0), .O(n121), .CO(n122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(208)
    defparam \tx_dac_fsm_inst/add_136/i2 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_136/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \fifo_inst/add_12/i2  (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[0] ), 
            .CI(1'b0), .O(n124), .CO(n125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \fifo_inst/add_12/i2 .I0_POLARITY = 1'b1;
    defparam \fifo_inst/add_12/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_fifo/add_12/i2  (.I0(\tx_fifo/wr_index[1] ), .I1(\tx_fifo/wr_index[0] ), 
            .CI(1'b0), .O(n147), .CO(n148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \tx_fifo/add_12/i2 .I0_POLARITY = 1'b1;
    defparam \tx_fifo/add_12/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \rx_fifo/add_12/i2  (.I0(\rx_fifo/wr_index[1] ), .I1(\rx_fifo/wr_index[0] ), 
            .CI(1'b0), .O(n193), .CO(n194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \rx_fifo/add_12/i2 .I0_POLARITY = 1'b1;
    defparam \rx_fifo/add_12/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \rx_fifo/add_12/i8  (.I0(\rx_fifo/wr_index[7] ), .I1(1'b0), 
            .CI(n3183), .O(n3179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \rx_fifo/add_12/i8 .I0_POLARITY = 1'b1;
    defparam \rx_fifo/add_12/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \rx_fifo/add_12/i7  (.I0(\rx_fifo/wr_index[6] ), .I1(1'b0), 
            .CI(n3186), .O(n3182), .CO(n3183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \rx_fifo/add_12/i7 .I0_POLARITY = 1'b1;
    defparam \rx_fifo/add_12/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \rx_fifo/add_12/i6  (.I0(\rx_fifo/wr_index[5] ), .I1(1'b0), 
            .CI(n3190), .O(n3185), .CO(n3186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \rx_fifo/add_12/i6 .I0_POLARITY = 1'b1;
    defparam \rx_fifo/add_12/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \rx_fifo/add_12/i5  (.I0(\rx_fifo/wr_index[4] ), .I1(1'b0), 
            .CI(n3193), .O(n3189), .CO(n3190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \rx_fifo/add_12/i5 .I0_POLARITY = 1'b1;
    defparam \rx_fifo/add_12/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \rx_fifo/add_12/i4  (.I0(\rx_fifo/wr_index[3] ), .I1(1'b0), 
            .CI(n3197), .O(n3192), .CO(n3193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \rx_fifo/add_12/i4 .I0_POLARITY = 1'b1;
    defparam \rx_fifo/add_12/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \rx_fifo/add_12/i3  (.I0(\rx_fifo/wr_index[2] ), .I1(1'b0), 
            .CI(n194), .O(n3196), .CO(n3197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \rx_fifo/add_12/i3 .I0_POLARITY = 1'b1;
    defparam \rx_fifo/add_12/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_fifo/add_12/i8  (.I0(\tx_fifo/wr_index[7] ), .I1(1'b0), 
            .CI(n3206), .O(n3202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \tx_fifo/add_12/i8 .I0_POLARITY = 1'b1;
    defparam \tx_fifo/add_12/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_fifo/add_12/i7  (.I0(\tx_fifo/wr_index[6] ), .I1(1'b0), 
            .CI(n3209), .O(n3205), .CO(n3206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \tx_fifo/add_12/i7 .I0_POLARITY = 1'b1;
    defparam \tx_fifo/add_12/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_fifo/add_12/i6  (.I0(\tx_fifo/wr_index[5] ), .I1(1'b0), 
            .CI(n3213), .O(n3208), .CO(n3209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \tx_fifo/add_12/i6 .I0_POLARITY = 1'b1;
    defparam \tx_fifo/add_12/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_fifo/add_12/i5  (.I0(\tx_fifo/wr_index[4] ), .I1(1'b0), 
            .CI(n3216), .O(n3212), .CO(n3213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \tx_fifo/add_12/i5 .I0_POLARITY = 1'b1;
    defparam \tx_fifo/add_12/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_fifo/add_12/i4  (.I0(\tx_fifo/wr_index[3] ), .I1(1'b0), 
            .CI(n3220), .O(n3215), .CO(n3216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \tx_fifo/add_12/i4 .I0_POLARITY = 1'b1;
    defparam \tx_fifo/add_12/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_fifo/add_12/i3  (.I0(\tx_fifo/wr_index[2] ), .I1(1'b0), 
            .CI(n148), .O(n3219), .CO(n3220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \tx_fifo/add_12/i3 .I0_POLARITY = 1'b1;
    defparam \tx_fifo/add_12/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \fifo_inst/add_12/i8  (.I0(\fifo_inst/wr_index[7] ), .I1(1'b0), 
            .CI(n3229), .O(n3226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \fifo_inst/add_12/i8 .I0_POLARITY = 1'b1;
    defparam \fifo_inst/add_12/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \fifo_inst/add_12/i7  (.I0(\fifo_inst/wr_index[6] ), .I1(1'b0), 
            .CI(n3232), .O(n3228), .CO(n3229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \fifo_inst/add_12/i7 .I0_POLARITY = 1'b1;
    defparam \fifo_inst/add_12/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \fifo_inst/add_12/i6  (.I0(\fifo_inst/wr_index[5] ), .I1(1'b0), 
            .CI(n3235), .O(n3231), .CO(n3232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \fifo_inst/add_12/i6 .I0_POLARITY = 1'b1;
    defparam \fifo_inst/add_12/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \fifo_inst/add_12/i5  (.I0(\fifo_inst/wr_index[4] ), .I1(1'b0), 
            .CI(n3238), .O(n3234), .CO(n3235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \fifo_inst/add_12/i5 .I0_POLARITY = 1'b1;
    defparam \fifo_inst/add_12/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \fifo_inst/add_12/i4  (.I0(\fifo_inst/wr_index[3] ), .I1(1'b0), 
            .CI(n3261), .O(n3237), .CO(n3238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \fifo_inst/add_12/i4 .I0_POLARITY = 1'b1;
    defparam \fifo_inst/add_12/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \fifo_inst/add_12/i3  (.I0(\fifo_inst/wr_index[2] ), .I1(1'b0), 
            .CI(n125), .O(n3260), .CO(n3261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\fifo.sv(51)
    defparam \fifo_inst/add_12/i3 .I0_POLARITY = 1'b1;
    defparam \fifo_inst/add_12/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_136/i6  (.I0(\tx_dac_fsm_inst/dctr[5] ), 
            .I1(1'b0), .CI(n3270), .O(n3267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(208)
    defparam \tx_dac_fsm_inst/add_136/i6 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_136/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_136/i5  (.I0(\tx_dac_fsm_inst/dctr[4] ), 
            .I1(1'b0), .CI(n3274), .O(n3269), .CO(n3270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(208)
    defparam \tx_dac_fsm_inst/add_136/i5 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_136/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_136/i4  (.I0(\tx_dac_fsm_inst/dctr[3] ), 
            .I1(1'b0), .CI(n7055), .O(n3273), .CO(n3274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(208)
    defparam \tx_dac_fsm_inst/add_136/i4 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_136/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_136/i3  (.I0(\tx_dac_fsm_inst/dctr[2] ), 
            .I1(1'b0), .CI(n122), .O(n3276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(208)
    defparam \tx_dac_fsm_inst/add_136/i3 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_136/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_129/i6  (.I0(\tx_dac_fsm_inst/zctr[5] ), 
            .I1(1'b0), .CI(n3285), .O(n3282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(197)
    defparam \tx_dac_fsm_inst/add_129/i6 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_129/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_129/i5  (.I0(\tx_dac_fsm_inst/zctr[4] ), 
            .I1(1'b0), .CI(n3289), .O(n3284), .CO(n3285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(197)
    defparam \tx_dac_fsm_inst/add_129/i5 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_129/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_129/i4  (.I0(\tx_dac_fsm_inst/zctr[3] ), 
            .I1(1'b0), .CI(n7056), .O(n3288), .CO(n3289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(197)
    defparam \tx_dac_fsm_inst/add_129/i4 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_129/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_129/i3  (.I0(\tx_dac_fsm_inst/zctr[2] ), 
            .I1(1'b0), .CI(n119), .O(n3295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(197)
    defparam \tx_dac_fsm_inst/add_129/i3 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_129/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/sub_20/add_2/i5  (.I0(\tx_dac_fsm_inst/sym_ctr[4] ), 
            .I1(1'b0), .CI(n7057), .O(n3300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(97)
    defparam \tx_dac_fsm_inst/sub_20/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sub_20/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/sub_20/add_2/i4  (.I0(\tx_dac_fsm_inst/sym_ctr[3] ), 
            .I1(1'b1), .CI(n7058), .O(n3302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(97)
    defparam \tx_dac_fsm_inst/sub_20/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/sub_20/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_18/i5  (.I0(\tx_dac_fsm_inst/sym_ctr[4] ), 
            .I1(1'b0), .CI(n3311), .O(n3307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(95)
    defparam \tx_dac_fsm_inst/add_18/i5 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_18/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_18/i4  (.I0(\tx_dac_fsm_inst/sym_ctr[3] ), 
            .I1(1'b0), .CI(n3314), .O(n3310), .CO(n3311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(95)
    defparam \tx_dac_fsm_inst/add_18/i4 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_18/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_18/i3  (.I0(\tx_dac_fsm_inst/sym_ctr[2] ), 
            .I1(1'b0), .CI(n3317), .O(n3313), .CO(n3314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(95)
    defparam \tx_dac_fsm_inst/add_18/i3 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_18/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \tx_dac_fsm_inst/add_18/i2  (.I0(\tx_dac_fsm_inst/sym_ctr[1] ), 
            .I1(1'b1), .CI(n7059), .O(n3316), .CO(n3317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(95)
    defparam \tx_dac_fsm_inst/add_18/i2 .I0_POLARITY = 1'b1;
    defparam \tx_dac_fsm_inst/add_18/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i24  (.I0(\led_inst/counter[23] ), .I1(1'b0), 
            .CI(n3327), .O(n3324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i24 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i23  (.I0(\led_inst/counter[22] ), .I1(1'b0), 
            .CI(n3330), .O(n3326), .CO(n3327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i23 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i22  (.I0(\led_inst/counter[21] ), .I1(1'b0), 
            .CI(n3334), .O(n3329), .CO(n3330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i22 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i21  (.I0(\led_inst/counter[20] ), .I1(1'b0), 
            .CI(n3340), .O(n3333), .CO(n3334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i21 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i20  (.I0(\led_inst/counter[19] ), .I1(1'b0), 
            .CI(n3344), .O(n3339), .CO(n3340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i20 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i19  (.I0(\led_inst/counter[18] ), .I1(1'b0), 
            .CI(n3347), .O(n3343), .CO(n3344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i19 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i18  (.I0(\led_inst/counter[17] ), .I1(1'b0), 
            .CI(n3351), .O(n3346), .CO(n3347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i18 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i17  (.I0(\led_inst/counter[16] ), .I1(1'b0), 
            .CI(n3358), .O(n3350), .CO(n3351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i17 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i16  (.I0(\led_inst/counter[15] ), .I1(1'b0), 
            .CI(n3363), .O(n3357), .CO(n3358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i16 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i15  (.I0(\led_inst/counter[14] ), .I1(1'b0), 
            .CI(n3367), .O(n3362), .CO(n3363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i15 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i14  (.I0(\led_inst/counter[13] ), .I1(1'b0), 
            .CI(n3371), .O(n3366), .CO(n3367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i14 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i13  (.I0(\led_inst/counter[12] ), .I1(1'b0), 
            .CI(n3376), .O(n3370), .CO(n3371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i13 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i12  (.I0(\led_inst/counter[11] ), .I1(1'b0), 
            .CI(n3380), .O(n3375), .CO(n3376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i12 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i11  (.I0(\led_inst/counter[10] ), .I1(1'b0), 
            .CI(n3386), .O(n3379), .CO(n3380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i11 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i10  (.I0(\led_inst/counter[9] ), .I1(1'b0), 
            .CI(n3390), .O(n3385), .CO(n3386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i10 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i9  (.I0(\led_inst/counter[8] ), .I1(1'b0), 
            .CI(n3393), .O(n3389), .CO(n3390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i9 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i8  (.I0(\led_inst/counter[7] ), .I1(1'b0), 
            .CI(n3397), .O(n3392), .CO(n3393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i8 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i7  (.I0(\led_inst/counter[6] ), .I1(1'b0), 
            .CI(n3400), .O(n3396), .CO(n3397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i7 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i6  (.I0(\led_inst/counter[5] ), .I1(1'b0), 
            .CI(n3404), .O(n3399), .CO(n3400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i6 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i5  (.I0(\led_inst/counter[4] ), .I1(1'b0), 
            .CI(n3407), .O(n3403), .CO(n3404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i5 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i4  (.I0(\led_inst/counter[3] ), .I1(1'b0), 
            .CI(n3411), .O(n3406), .CO(n3407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i4 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \led_inst/add_23/i3  (.I0(\led_inst/counter[2] ), .I1(1'b0), 
            .CI(n20), .O(n3410), .CO(n3411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\led.sv(78)
    defparam \led_inst/add_23/i3 .I0_POLARITY = 1'b1;
    defparam \led_inst/add_23/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \spi_slave_inst/add_29/i5  (.I0(\spi_slave_inst/bitcnt[4] ), .I1(1'b0), 
            .CI(n3420), .O(n3416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/add_29/i5 .I0_POLARITY = 1'b1;
    defparam \spi_slave_inst/add_29/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \spi_slave_inst/add_29/i4  (.I0(\spi_slave_inst/bitcnt[3] ), .I1(1'b0), 
            .CI(n3423), .O(n3419), .CO(n3420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/add_29/i4 .I0_POLARITY = 1'b1;
    defparam \spi_slave_inst/add_29/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \spi_slave_inst/add_29/i3  (.I0(\spi_slave_inst/bitcnt[2] ), .I1(1'b0), 
            .CI(n3427), .O(n3422), .CO(n3423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/add_29/i3 .I0_POLARITY = 1'b1;
    defparam \spi_slave_inst/add_29/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \spi_slave_inst/add_29/i2  (.I0(\spi_slave_inst/bitcnt[1] ), .I1(\spi_slave_inst/bitcnt[0] ), 
            .CI(1'b0), .O(n3426), .CO(n3427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\spi_slave.sv(92)
    defparam \spi_slave_inst/add_29/i2 .I0_POLARITY = 1'b1;
    defparam \spi_slave_inst/add_29/i2 .I1_POLARITY = 1'b1;
    EFX_LUT4 LUT__7664 (.I0(\gpo_inst/gp_config_reg[6] ), .I1(\gpo_inst/gp_config_reg[7] ), 
            .O(gpo_pins[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7664.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7665 (.I0(\gpo_inst/gp_config_reg[5] ), .I1(\gpo_inst/gp_config_reg[7] ), 
            .O(gpo_pins[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7665.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7666 (.I0(\gpo_inst/gp_config_reg[4] ), .I1(\gpo_inst/gp_config_reg[7] ), 
            .O(gpo_pins[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7666.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7667 (.I0(\gpo_inst/gp_config_reg[3] ), .I1(\gpo_inst/gp_config_reg[7] ), 
            .O(gpo_pins[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7667.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7668 (.I0(\gpo_inst/gp_config_reg[2] ), .I1(\gpo_inst/gp_config_reg[7] ), 
            .O(gpo_pins[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7668.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7669 (.I0(\gpo_inst/gp_config_reg[1] ), .I1(\gpo_inst/gp_config_reg[7] ), 
            .O(gpo_pins[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7669.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7670 (.I0(\gpo_inst/gp_config_reg[0] ), .I1(\gpo_inst/gp_config_reg[7] ), 
            .O(gpo_pins[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7670.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7671 (.I0(\tx_dac_fsm_inst/dac_config_reg[0] ), .I1(n136), 
            .O(lvds_tx_inst1_DATA[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7671.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7672 (.I0(n116), .I1(\tx_dac_fsm_inst/dac_config_reg[0] ), 
            .O(lvds_tx_inst1_DATA[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7672.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7673 (.I0(\spi_slave_inst/sync_ss[1] ), .I1(\spi_slave_inst/sync_ss[2] ), 
            .O(n4236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7673.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7674 (.I0(n4236), .I1(\reg_addr[3] ), .O(\spi_slave_inst/n94 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7674.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7675 (.I0(\spi_slave_inst/bitcnt[2] ), .I1(\spi_slave_inst/bitcnt[1] ), 
            .I2(\spi_slave_inst/bitcnt[0] ), .O(n4237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__7675.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__7676 (.I0(\spi_slave_inst/sync_sclk[2] ), .I1(\spi_slave_inst/sync_ss[1] ), 
            .I2(\spi_slave_inst/sync_sclk[1] ), .O(n4238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7676.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7677 (.I0(n4237), .I1(n4238), .I2(n4235), .I3(n4236), 
            .O(ceg_net49)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__7677.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__7678 (.I0(n4236), .I1(\reg_addr[2] ), .O(\spi_slave_inst/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7678.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7679 (.I0(n4236), .I1(n3422), .O(\spi_slave_inst/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7679.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7680 (.I0(n4236), .I1(n4238), .O(ceg_net40)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7680.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7681 (.I0(n4236), .I1(n3426), .O(\spi_slave_inst/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7681.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7682 (.I0(n4236), .I1(\reg_addr[1] ), .O(\spi_slave_inst/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7682.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7683 (.I0(n4236), .I1(\reg_addr[0] ), .O(\spi_slave_inst/n97 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7683.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7684 (.I0(\reg_addr[4] ), .I1(\reg_addr[3] ), .I2(\reg_addr[5] ), 
            .I3(\reg_addr[6] ), .O(n4239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__7684.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__7685 (.I0(\reg_addr[2] ), .I1(\reg_addr[1] ), .I2(\reg_addr[5] ), 
            .I3(\reg_addr[6] ), .O(n4240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__7685.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__7686 (.I0(\reg_addr[4] ), .I1(n4240), .I2(\reg_addr[3] ), 
            .O(n4241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__7686.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__7687 (.I0(rw_out), .I1(addr_dv), .O(n4242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7687.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7688 (.I0(n4241), .I1(n4239), .I2(n4242), .O(tx_en)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__7688.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__7689 (.I0(n4236), .I1(\spi_slave_inst/bitcnt[0] ), .O(\spi_slave_inst/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7689.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7690 (.I0(\spi_slave_inst/sync_ss[1] ), .I1(\spi_slave_inst/sync_ss[2] ), 
            .O(\spi_slave_inst/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__7690.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__7691 (.I0(\spi_slave_inst/n68 ), .I1(\spi_slave_inst/sync_mosi[1] ), 
            .O(\spi_slave_inst/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7691.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7692 (.I0(n4238), .I1(n4235), .I2(n4237), .I3(\spi_slave_inst/n68 ), 
            .O(ceg_net23)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__7692.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__7693 (.I0(n4236), .I1(\spi_slave_inst/sync_mosi[1] ), 
            .O(\spi_slave_inst/n98 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7693.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7694 (.I0(\reg_addr[0] ), .I1(n4242), .O(n4243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7694.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7695 (.I0(\reg_addr[2] ), .I1(\reg_addr[1] ), .I2(n4243), 
            .I3(n4239), .O(n4244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__7695.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__7696 (.I0(\reg_addr[2] ), .I1(n4239), .I2(n4242), .I3(\reg_addr[1] ), 
            .O(n4245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__7696.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__7697 (.I0(\tx_fifo/buff_head[0] ), .I1(\reg_addr[0] ), 
            .I2(n4245), .O(n4246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__7697.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__7698 (.I0(\reg_addr[1] ), .I1(\reg_addr[2] ), .O(n4247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7698.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7699 (.I0(n4239), .I1(n4247), .O(n4248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7699.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7700 (.I0(\rx_fifo/length[0] ), .I1(\rx_fifo/buff_head[0] ), 
            .I2(\reg_addr[0] ), .I3(n4248), .O(n4249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__7700.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__7701 (.I0(\fifo_inst/length[0] ), .I1(\fifo_inst/buff_head[0] ), 
            .I2(\reg_addr[0] ), .I3(n4241), .O(n4250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__7701.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__7702 (.I0(n4239), .I1(\reg_addr[2] ), .I2(\reg_addr[1] ), 
            .O(n4251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__7702.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__7703 (.I0(\tx_dac_fsm_inst/dac_config_reg[0] ), .I1(\data_from_led[0] ), 
            .I2(\reg_addr[0] ), .I3(n4251), .O(n4252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__7703.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__7704 (.I0(n4249), .I1(n4250), .I2(n4252), .I3(n4242), 
            .O(n4253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__7704.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__7705 (.I0(\reg_addr[2] ), .I1(\tx_fifo/length[0] ), .I2(\reg_addr[1] ), 
            .I3(n4243), .O(n4254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__7705.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__7706 (.I0(n4253), .I1(n4246), .I2(n4254), .O(n4255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__7706.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__7707 (.I0(\spi_slave_inst/sync_tx_en[1] ), .I1(\spi_slave_inst/sync_tx_en[0] ), 
            .O(n4256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7707.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7708 (.I0(\gpo_inst/gp_config_reg[0] ), .I1(n4244), .I2(n4255), 
            .I3(n4256), .O(\spi_slave_inst/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__7708.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__7709 (.I0(n4238), .I1(n4256), .I2(tx_en), .O(ceg_net77)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7709.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7710 (.I0(rw_out), .I1(n4235), .I2(n4238), .I3(n4236), 
            .O(ceg_net98)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__7710.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__7711 (.I0(\spi_slave_inst/n68 ), .I1(n4235), .O(ceg_net34)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7711.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7712 (.I0(\spi_slave_inst/sync_sclk[2] ), .I1(\spi_slave_inst/bitcnt[1] ), 
            .I2(\spi_slave_inst/sync_sclk[1] ), .I3(\spi_slave_inst/bitcnt[2] ), 
            .O(n4257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__7712.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__7713 (.I0(rw_out), .I1(\spi_slave_inst/bitcnt[4] ), .I2(\spi_slave_inst/bitcnt[0] ), 
            .I3(\spi_slave_inst/bitcnt[3] ), .O(n4258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__7713.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__7714 (.I0(n4258), .I1(n4257), .I2(\spi_slave_inst/n68 ), 
            .O(ceg_net37)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__7714.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__7715 (.I0(n4236), .I1(n3416), .O(\spi_slave_inst/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7715.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7716 (.I0(n4236), .I1(\reg_addr[4] ), .O(\spi_slave_inst/n93 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7716.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7717 (.I0(n4236), .I1(n3419), .O(\spi_slave_inst/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7717.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7718 (.I0(n4236), .I1(\reg_addr[5] ), .O(\spi_slave_inst/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7718.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7719 (.I0(n4256), .I1(n4238), .I2(tx_en), .O(n4259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__7719.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__7720 (.I0(\tx_fifo/length[1] ), .I1(\tx_fifo/buff_head[1] ), 
            .I2(\reg_addr[0] ), .I3(n4245), .O(n4260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__7720.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__7721 (.I0(\reg_addr[2] ), .I1(\rx_fifo/length[1] ), .I2(\reg_addr[1] ), 
            .I3(n4239), .O(n4261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__7721.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__7722 (.I0(\rx_fifo/buff_head[1] ), .I1(n4248), .I2(n4261), 
            .I3(\reg_addr[0] ), .O(n4262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__7722.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__7723 (.I0(n4243), .I1(n4251), .O(n4263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7723.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7724 (.I0(n4262), .I1(n4242), .I2(\data_from_led[1] ), 
            .I3(n4263), .O(n4264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__7724.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__7725 (.I0(n4241), .I1(n4242), .O(n4265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7725.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7726 (.I0(\fifo_inst/length[1] ), .I1(\fifo_inst/buff_head[1] ), 
            .I2(\reg_addr[0] ), .I3(n4265), .O(n4266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__7726.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__7727 (.I0(n4244), .I1(\gpo_inst/gp_config_reg[1] ), .I2(n4256), 
            .O(n4267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7727.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7728 (.I0(n4266), .I1(n4260), .I2(n4264), .I3(n4267), 
            .O(n4268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__7728.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__7729 (.I0(\spi_slave_inst/d_o[0] ), .I1(n4259), .I2(n4268), 
            .O(\spi_slave_inst/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8 */ ;
    defparam LUT__7729.LUTMASK = 16'hf8f8;
    EFX_LUT4 LUT__7730 (.I0(n4248), .I1(n4242), .I2(\reg_addr[0] ), .O(n4269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__7730.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__7731 (.I0(n4243), .I1(n4248), .O(n4270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7731.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7732 (.I0(n4270), .I1(\rx_fifo/length[2] ), .I2(n4269), 
            .I3(\rx_fifo/buff_head[2] ), .O(n4271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__7732.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__7733 (.I0(n4263), .I1(\data_from_led[2] ), .I2(n4271), 
            .O(n4272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__7733.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__7734 (.I0(\tx_fifo/buff_head[2] ), .I1(\tx_fifo/length[2] ), 
            .I2(\reg_addr[0] ), .I3(n4245), .O(n4273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__7734.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__7735 (.I0(\fifo_inst/length[2] ), .I1(\fifo_inst/buff_head[2] ), 
            .I2(\reg_addr[0] ), .I3(n4265), .O(n4274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__7735.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__7736 (.I0(n4244), .I1(\gpo_inst/gp_config_reg[2] ), .I2(n4273), 
            .I3(n4274), .O(n4275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__7736.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__7737 (.I0(n4259), .I1(\spi_slave_inst/d_o[1] ), .O(n4276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7737.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7738 (.I0(n4275), .I1(n4272), .I2(n4256), .I3(n4276), 
            .O(\spi_slave_inst/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff70 */ ;
    defparam LUT__7738.LUTMASK = 16'hff70;
    EFX_LUT4 LUT__7739 (.I0(\tx_fifo/length[3] ), .I1(\tx_fifo/buff_head[3] ), 
            .I2(\reg_addr[0] ), .I3(n4245), .O(n4277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__7739.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__7740 (.I0(\reg_addr[2] ), .I1(\rx_fifo/length[3] ), .I2(\reg_addr[1] ), 
            .I3(n4239), .O(n4278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__7740.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__7741 (.I0(\rx_fifo/buff_head[3] ), .I1(n4248), .I2(n4278), 
            .I3(\reg_addr[0] ), .O(n4279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__7741.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__7742 (.I0(n4279), .I1(n4242), .I2(\data_from_led[3] ), 
            .I3(n4263), .O(n4280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__7742.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__7743 (.I0(\fifo_inst/length[3] ), .I1(\fifo_inst/buff_head[3] ), 
            .I2(\reg_addr[0] ), .I3(n4265), .O(n4281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__7743.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__7744 (.I0(n4244), .I1(\gpo_inst/gp_config_reg[3] ), .I2(n4256), 
            .O(n4282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7744.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7745 (.I0(n4281), .I1(n4277), .I2(n4280), .I3(n4282), 
            .O(n4283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__7745.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__7746 (.I0(\spi_slave_inst/d_o[2] ), .I1(n4259), .I2(n4283), 
            .O(\spi_slave_inst/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8 */ ;
    defparam LUT__7746.LUTMASK = 16'hf8f8;
    EFX_LUT4 LUT__7747 (.I0(\reg_addr[2] ), .I1(\rx_fifo/length[4] ), .I2(\reg_addr[1] ), 
            .I3(n4239), .O(n4284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__7747.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__7748 (.I0(\rx_fifo/buff_head[4] ), .I1(n4248), .I2(n4284), 
            .I3(\reg_addr[0] ), .O(n4285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__7748.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__7749 (.I0(\fifo_inst/length[4] ), .I1(\fifo_inst/buff_head[4] ), 
            .I2(\reg_addr[0] ), .I3(n4265), .O(n4286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__7749.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__7750 (.I0(\tx_fifo/buff_head[4] ), .I1(\tx_fifo/length[4] ), 
            .I2(\reg_addr[0] ), .O(n4287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7750.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7751 (.I0(n4263), .I1(\data_from_led[4] ), .I2(n4287), 
            .I3(n4245), .O(n4288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__7751.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__7752 (.I0(n4285), .I1(n4242), .I2(n4286), .I3(n4288), 
            .O(n4289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__7752.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__7753 (.I0(n4244), .I1(\gpo_inst/gp_config_reg[4] ), .I2(n4256), 
            .O(n4290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__7753.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__7754 (.I0(n4289), .I1(n4290), .I2(n4259), .I3(\spi_slave_inst/d_o[3] ), 
            .O(\spi_slave_inst/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__7754.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__7755 (.I0(\tx_fifo/buff_head[5] ), .I1(\tx_fifo/length[5] ), 
            .I2(\reg_addr[0] ), .I3(n4245), .O(n4291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__7755.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__7756 (.I0(n4263), .I1(\data_from_led[5] ), .I2(n4291), 
            .O(n4292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__7756.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__7757 (.I0(n4270), .I1(\rx_fifo/length[5] ), .I2(n4269), 
            .I3(\rx_fifo/buff_head[5] ), .O(n4293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__7757.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__7758 (.I0(\fifo_inst/length[5] ), .I1(\fifo_inst/buff_head[5] ), 
            .I2(\reg_addr[0] ), .O(n4294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7758.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7759 (.I0(n4294), .I1(n4265), .I2(n4244), .I3(\gpo_inst/gp_config_reg[5] ), 
            .O(n4295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__7759.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__7760 (.I0(n4293), .I1(n4295), .I2(n4292), .I3(n4256), 
            .O(n4296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__7760.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__7761 (.I0(\spi_slave_inst/d_o[4] ), .I1(n4259), .I2(n4296), 
            .O(\spi_slave_inst/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8 */ ;
    defparam LUT__7761.LUTMASK = 16'hf8f8;
    EFX_LUT4 LUT__7762 (.I0(\fifo_inst/length[6] ), .I1(\fifo_inst/buff_head[6] ), 
            .I2(\reg_addr[0] ), .I3(n4265), .O(n4297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__7762.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__7764 (.I0(n4263), .I1(n4269), .O(n4298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7764.LUTMASK = 16'h1111;
    EFX_LUT4 \tx_dac_fsm_inst/dlatchrs_162/i1  (.I0(n3556), .I1(n109), .I2(n3557), 
            .O(n109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam \tx_dac_fsm_inst/dlatchrs_162/i1 .LUTMASK = 16'hacac;
    EFX_LUT4 LUT__7765 (.I0(\data_from_led[6] ), .I1(n4263), .I2(\rx_fifo/buff_head[6] ), 
            .I3(n4269), .O(n4299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__7765.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__7766 (.I0(n4243), .I1(n4248), .I2(\rx_fifo/length[6] ), 
            .O(n4300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__7766.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__7767 (.I0(\tx_fifo/buff_head[6] ), .I1(\tx_fifo/length[6] ), 
            .I2(\reg_addr[0] ), .I3(n4245), .O(n4301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__7767.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__7768 (.I0(n4244), .I1(\gpo_inst/gp_config_reg[6] ), .I2(n4300), 
            .I3(n4301), .O(n4302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__7768.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__7769 (.I0(n4297), .I1(n4298), .I2(n4299), .I3(n4302), 
            .O(n4303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__7769.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__7770 (.I0(n4303), .I1(n4256), .I2(n4259), .I3(\spi_slave_inst/d_o[5] ), 
            .O(\spi_slave_inst/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__7770.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__7771 (.I0(\fifo_inst/length[7] ), .I1(\fifo_inst/buff_head[7] ), 
            .I2(\reg_addr[0] ), .I3(n4265), .O(n4304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__7771.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__7772 (.I0(\data_from_led[7] ), .I1(n4263), .I2(\rx_fifo/buff_head[7] ), 
            .I3(n4269), .O(n4305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__7772.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__7773 (.I0(n4243), .I1(n4248), .I2(\rx_fifo/length[7] ), 
            .O(n4306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__7773.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__7774 (.I0(\tx_fifo/buff_head[7] ), .I1(\tx_fifo/length[7] ), 
            .I2(\reg_addr[0] ), .I3(n4245), .O(n4307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__7774.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__7775 (.I0(n4244), .I1(\gpo_inst/gp_config_reg[7] ), .I2(n4306), 
            .I3(n4307), .O(n4308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__7775.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__7776 (.I0(n4304), .I1(n4298), .I2(n4305), .I3(n4308), 
            .O(n4309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__7776.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__7777 (.I0(n4309), .I1(n4256), .I2(n4259), .I3(\spi_slave_inst/d_o[6] ), 
            .O(\spi_slave_inst/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__7777.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__7778 (.I0(n4236), .I1(\rx_d[0] ), .O(\spi_slave_inst/n173 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7778.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7779 (.I0(n4236), .I1(\rx_d[1] ), .O(\spi_slave_inst/n172 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7779.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7780 (.I0(n4236), .I1(\rx_d[2] ), .O(\spi_slave_inst/n171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7780.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7781 (.I0(n4236), .I1(\rx_d[3] ), .O(\spi_slave_inst/n170 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7781.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7782 (.I0(n4236), .I1(\rx_d[4] ), .O(\spi_slave_inst/n169 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7782.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7783 (.I0(n4236), .I1(\rx_d[5] ), .O(\spi_slave_inst/n168 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7783.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7784 (.I0(n4236), .I1(\rx_d[6] ), .O(\spi_slave_inst/n167 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7784.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7785 (.I0(n4263), .I1(\led_inst/ctr_cfg_reg[7] ), .O(\led_inst/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7785.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7786 (.I0(n4263), .I1(\led_inst/ctr_cfg_reg[6] ), .O(\led_inst/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7786.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7787 (.I0(n4263), .I1(\led_inst/ctr_cfg_reg[5] ), .O(\led_inst/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7787.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7788 (.I0(n4263), .I1(\led_inst/ctr_cfg_reg[4] ), .O(\led_inst/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7788.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7789 (.I0(n4263), .I1(\led_inst/ctr_cfg_reg[3] ), .O(\led_inst/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7789.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7790 (.I0(n4263), .I1(\led_inst/ctr_cfg_reg[0] ), .O(\led_inst/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7790.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7791 (.I0(n4263), .I1(\led_inst/ctr_cfg_reg[2] ), .O(\led_inst/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7791.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7792 (.I0(n4263), .I1(\led_inst/ctr_cfg_reg[1] ), .O(\led_inst/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7792.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7793 (.I0(\led_inst/counter[17] ), .I1(\led_inst/counter[16] ), 
            .I2(\led_inst/ctr_cfg_reg[1] ), .I3(\led_inst/ctr_cfg_reg[0] ), 
            .O(n4310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__7793.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__7794 (.I0(\led_inst/counter[19] ), .I1(\led_inst/ctr_cfg_reg[3] ), 
            .O(n4311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7794.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7795 (.I0(n4310), .I1(\led_inst/ctr_cfg_reg[2] ), .I2(\led_inst/counter[18] ), 
            .I3(n4311), .O(n4312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__7795.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__7796 (.I0(\led_inst/ctr_cfg_reg[3] ), .I1(\led_inst/counter[19] ), 
            .I2(\led_inst/ctr_cfg_reg[4] ), .I3(\led_inst/counter[20] ), 
            .O(n4313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__7796.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__7797 (.I0(\led_inst/counter[20] ), .I1(\led_inst/ctr_cfg_reg[4] ), 
            .I2(\led_inst/counter[21] ), .I3(\led_inst/ctr_cfg_reg[5] ), 
            .O(n4314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__7797.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__7798 (.I0(\led_inst/ctr_cfg_reg[5] ), .I1(\led_inst/counter[21] ), 
            .I2(\led_inst/ctr_cfg_reg[6] ), .I3(\led_inst/counter[22] ), 
            .O(n4315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__7798.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__7799 (.I0(n4312), .I1(n4313), .I2(n4314), .I3(n4315), 
            .O(n4316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__7799.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__7800 (.I0(\led_inst/counter[22] ), .I1(\led_inst/ctr_cfg_reg[6] ), 
            .I2(n4316), .O(n4317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__7800.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__7801 (.I0(n4317), .I1(\led_inst/ctr_cfg_reg[7] ), .I2(\led_inst/counter[23] ), 
            .O(\led_inst/LessThan_21/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__7801.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__7802 (.I0(\led_inst/LessThan_21/n48 ), .I1(\led_inst/counter[0] ), 
            .O(\led_inst/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7802.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7803 (.I0(rw_out), .I1(\reg_addr[0] ), .I2(addr_dv), 
            .I3(rxdv), .O(n4318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__7803.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__7804 (.I0(n4251), .I1(n4318), .O(rx_en_led)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7804.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7805 (.I0(rx_en_led), .I1(\rx_d[0] ), .O(\data_to_led[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7805.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7806 (.I0(\led_inst/LessThan_21/n48 ), .I1(n19), .O(\led_inst/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7806.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7807 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3410), .O(\led_inst/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7807.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7808 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3406), .O(\led_inst/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7808.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7809 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3403), .O(\led_inst/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7809.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7810 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3399), .O(\led_inst/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7810.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7811 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3396), .O(\led_inst/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7811.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7812 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3392), .O(\led_inst/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7812.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7813 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3389), .O(\led_inst/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7813.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7814 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3385), .O(\led_inst/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7814.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7815 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3379), .O(\led_inst/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7815.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7816 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3375), .O(\led_inst/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7816.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7817 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3370), .O(\led_inst/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7817.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7818 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3366), .O(\led_inst/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7818.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7819 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3362), .O(\led_inst/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7819.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7820 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3357), .O(\led_inst/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7820.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7821 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3350), .O(\led_inst/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7821.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7822 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3346), .O(\led_inst/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7822.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7823 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3343), .O(\led_inst/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7823.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7824 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3339), .O(\led_inst/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7824.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7825 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3333), .O(\led_inst/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7825.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7826 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3329), .O(\led_inst/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7826.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7827 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3326), .O(\led_inst/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7827.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7828 (.I0(\led_inst/LessThan_21/n48 ), .I1(n3324), .O(\led_inst/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7828.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7829 (.I0(rx_en_led), .I1(\rx_d[1] ), .O(\data_to_led[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7829.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7830 (.I0(rx_en_led), .I1(\rx_d[2] ), .O(\data_to_led[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7830.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7831 (.I0(rx_en_led), .I1(\rx_d[3] ), .O(\data_to_led[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7831.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7832 (.I0(rx_en_led), .I1(\rx_d[4] ), .O(\data_to_led[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7832.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7833 (.I0(rx_en_led), .I1(\rx_d[5] ), .O(\data_to_led[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7833.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7834 (.I0(rx_en_led), .I1(\rx_d[6] ), .O(\data_to_led[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7834.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7835 (.I0(rx_en_led), .I1(\rx_d[7] ), .O(\data_to_led[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7835.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7836 (.I0(\reg_addr[2] ), .I1(\reg_addr[1] ), .I2(n4239), 
            .I3(n4318), .O(rx_en_gpo)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__7836.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__7837 (.I0(rx_en_gpo), .I1(\rx_d[0] ), .O(\data_to_gpo[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7837.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7838 (.I0(rx_en_gpo), .I1(\rx_d[1] ), .O(\data_to_gpo[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7838.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7839 (.I0(rx_en_gpo), .I1(\rx_d[2] ), .O(\data_to_gpo[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7839.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7840 (.I0(rx_en_gpo), .I1(\rx_d[3] ), .O(\data_to_gpo[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7840.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7841 (.I0(rx_en_gpo), .I1(\rx_d[4] ), .O(\data_to_gpo[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7841.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7842 (.I0(rx_en_gpo), .I1(\rx_d[5] ), .O(\data_to_gpo[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7842.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7843 (.I0(rx_en_gpo), .I1(\rx_d[6] ), .O(\data_to_gpo[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7843.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7844 (.I0(rx_en_gpo), .I1(\rx_d[7] ), .O(\data_to_gpo[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7844.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7845 (.I0(n4241), .I1(n4318), .O(rx_en_fifo)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7845.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7846 (.I0(rx_en_fifo), .I1(\rx_d[2] ), .O(\data_to_fifo[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7846.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7847 (.I0(\fifo_inst/sync_wr[1] ), .I1(\fifo_inst/sync_wr[0] ), 
            .O(n4319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7847.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7848 (.I0(\fifo_inst/wr_index[7] ), .I1(\fifo_inst/wr_index[0] ), 
            .I2(n4319), .O(n4320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__7848.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__7849 (.I0(\fifo_inst/wr_index[5] ), .I1(\fifo_inst/wr_index[6] ), 
            .I2(n4320), .O(n4321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7849.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7850 (.I0(\fifo_inst/wr_index[2] ), .I1(\fifo_inst/wr_index[3] ), 
            .I2(\fifo_inst/wr_index[4] ), .I3(\fifo_inst/wr_index[1] ), 
            .O(n4322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__7850.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__7851 (.I0(n4321), .I1(n4322), .O(\i14/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7851.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7852 (.I0(rx_en_fifo), .I1(\rx_d[1] ), .O(\data_to_fifo[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7852.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7853 (.I0(rx_en_fifo), .I1(\rx_d[0] ), .O(\data_to_fifo[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7853.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7854 (.I0(rx_en_fifo), .I1(\rx_d[7] ), .O(\data_to_fifo[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7854.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7855 (.I0(\fifo_inst/wr_index[0] ), .I1(\fifo_inst/wr_index[7] ), 
            .I2(n4319), .O(n4323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7855.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7856 (.I0(\fifo_inst/wr_index[5] ), .I1(\fifo_inst/wr_index[6] ), 
            .I2(n4323), .O(n4324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7856.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7857 (.I0(n4324), .I1(n4322), .O(\i14/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7857.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7858 (.I0(\tx_dac_fsm_inst/sym_ctr[2] ), .I1(\tx_dac_fsm_inst/sym_ctr[3] ), 
            .O(n4167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__7858.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__7859 (.I0(n4167), .I1(\tx_dac_fsm_inst/sym_ctr[4] ), .O(n4325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7859.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7860 (.I0(n4325), .I1(\tx_dac_fsm_inst/sym_ctr[0] ), .O(\tx_dac_fsm_inst/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__7860.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__7861 (.I0(\tx_dac_fsm_inst/zctr[0] ), .I1(\tx_dac_fsm_inst/zctr[1] ), 
            .I2(\tx_dac_fsm_inst/zctr[2] ), .O(n4161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__7861.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__7862 (.I0(\tx_dac_fsm_inst/zctr[4] ), .I1(\tx_dac_fsm_inst/zctr[5] ), 
            .I2(n4161), .I3(\tx_dac_fsm_inst/zctr[3] ), .O(n4326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__7862.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__7863 (.I0(\tx_dac_fsm_inst/dctr[1] ), .I1(\tx_dac_fsm_inst/dctr[2] ), 
            .O(n4327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7863.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7864 (.I0(n4327), .I1(\tx_dac_fsm_inst/dctr[0] ), .O(n4152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7864.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7865 (.I0(\tx_dac_fsm_inst/dctr[4] ), .I1(\tx_dac_fsm_inst/dctr[5] ), 
            .O(n4328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7865.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7866 (.I0(n4152), .I1(n4328), .I2(\tx_dac_fsm_inst/dctr[3] ), 
            .O(n4329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__7866.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__7867 (.I0(n4329), .I1(n4326), .I2(\tx_dac_fsm_inst/dac_config_reg[0] ), 
            .O(\tx_dac_fsm_inst/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__7867.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__7868 (.I0(\tx_dac_fsm_inst/n42 ), .I1(n4325), .O(\tx_dac_fsm_inst/n344 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7868.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7869 (.I0(\tx_dac_fsm_inst/sym_pos[2] ), .I1(\tx_dac_fsm_inst/sym_pos[1] ), 
            .I2(\tx_dac_fsm_inst/sym_pos[3] ), .I3(\tx_dac_fsm_inst/sym_pos[0] ), 
            .O(n4330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcf15 */ ;
    defparam LUT__7869.LUTMASK = 16'hcf15;
    EFX_LUT4 LUT__7870 (.I0(n4330), .I1(\tx_dac_fsm_inst/dac_config_reg[0] ), 
            .I2(\tx_dac_fsm_inst/state_reg[0] ), .I3(\tx_dac_fsm_inst/state_reg[1] ), 
            .O(n4331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__7870.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__7871 (.I0(\tx_dac_fsm_inst/dctr[3] ), .I1(n4327), .I2(n4328), 
            .I3(\tx_dac_fsm_inst/state_reg[0] ), .O(n4332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__7871.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__7872 (.I0(n4332), .I1(\tx_dac_fsm_inst/state_reg[0] ), 
            .I2(\tx_dac_fsm_inst/state_reg[2] ), .I3(\tx_dac_fsm_inst/state_reg[3] ), 
            .O(n4333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfa3f */ ;
    defparam LUT__7872.LUTMASK = 16'hfa3f;
    EFX_LUT4 LUT__7873 (.I0(n4327), .I1(\tx_dac_fsm_inst/dctr[3] ), .I2(n4328), 
            .O(n4334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7873.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7874 (.I0(\tx_dac_fsm_inst/dctr[0] ), .I1(\tx_dac_fsm_inst/dctr[2] ), 
            .I2(\tx_dac_fsm_inst/state_reg[2] ), .I3(n4334), .O(n4335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__7874.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__7875 (.I0(\tx_dac_fsm_inst/state_reg[2] ), .I1(\tx_dac_fsm_inst/zctr[4] ), 
            .I2(\tx_dac_fsm_inst/zctr[5] ), .O(n4336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__7875.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__7876 (.I0(\tx_dac_fsm_inst/dac_config_reg[0] ), .I1(\tx_dac_fsm_inst/state_reg[2] ), 
            .O(n4337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7876.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7877 (.I0(\tx_dac_fsm_inst/state_reg[0] ), .I1(n4335), 
            .I2(n4336), .I3(n4337), .O(n4338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f1 */ ;
    defparam LUT__7877.LUTMASK = 16'h00f1;
    EFX_LUT4 LUT__7878 (.I0(n4338), .I1(n4333), .I2(\tx_dac_fsm_inst/state_reg[1] ), 
            .I3(\tx_dac_fsm_inst/state_reg[3] ), .O(n4339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc05 */ ;
    defparam LUT__7878.LUTMASK = 16'hfc05;
    EFX_LUT4 LUT__7879 (.I0(n4331), .I1(\tx_dac_fsm_inst/state_reg[2] ), 
            .I2(n4339), .O(n3556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__7879.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__7880 (.I0(\tx_dac_fsm_inst/state_reg[0] ), .I1(n4334), 
            .I2(\tx_dac_fsm_inst/state_reg[1] ), .I3(\tx_dac_fsm_inst/state_reg[2] ), 
            .O(n4340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__7880.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__7881 (.I0(n4337), .I1(\tx_dac_fsm_inst/state_reg[0] ), 
            .I2(\tx_dac_fsm_inst/state_reg[1] ), .I3(\tx_dac_fsm_inst/state_reg[3] ), 
            .O(n4341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__7881.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__7882 (.I0(n4340), .I1(n4341), .O(n3557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__7882.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__7883 (.I0(\tx_dac_fsm_inst/sym_ctr[1] ), .I1(n3316), .I2(n4325), 
            .O(\tx_dac_fsm_inst/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__7883.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__7884 (.I0(\tx_dac_fsm_inst/sym_ctr[2] ), .I1(n3313), .I2(n4325), 
            .O(\tx_dac_fsm_inst/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__7884.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__7885 (.I0(n3302), .I1(n3310), .I2(n4325), .O(\tx_dac_fsm_inst/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__7885.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__7886 (.I0(\tx_dac_fsm_inst/state_reg[0] ), .I1(\tx_dac_fsm_inst/state_reg[1] ), 
            .I2(\tx_dac_fsm_inst/state_reg[2] ), .I3(\tx_dac_fsm_inst/state_reg[3] ), 
            .O(n3561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__7886.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__7887 (.I0(\tx_dac_fsm_inst/state_reg[1] ), .I1(\tx_dac_fsm_inst/state_reg[2] ), 
            .O(n4342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7887.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7888 (.I0(n4342), .I1(\tx_dac_fsm_inst/state_reg[3] ), 
            .O(n3562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__7888.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__7889 (.I0(rx_en_fifo), .I1(\rx_d[6] ), .O(\data_to_fifo[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7889.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7890 (.I0(\tx_dac_fsm_inst/state_reg[3] ), .I1(\tx_dac_fsm_inst/state_reg[0] ), 
            .I2(n4342), .O(n3564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__7890.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__7891 (.I0(\tx_dac_fsm_inst/state_reg[2] ), .I1(\tx_dac_fsm_inst/state_reg[1] ), 
            .I2(\tx_dac_fsm_inst/state_reg[0] ), .O(n3565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__7891.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__7892 (.I0(\tx_dac_fsm_inst/zctr[0] ), .I1(n115), .O(\tx_dac_fsm_inst/n258 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7892.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7893 (.I0(n3300), .I1(n3307), .I2(n4325), .O(\tx_dac_fsm_inst/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__7893.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__7894 (.I0(\tx_dac_fsm_inst/dctr[0] ), .I1(n113), .O(\tx_dac_fsm_inst/n284 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7894.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7895 (.I0(rw_out), .I1(\reg_addr[0] ), .I2(addr_dv), 
            .I3(rxdv), .O(n4343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__7895.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__7896 (.I0(n4251), .I1(n4343), .O(rx_en_dac)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7896.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7897 (.I0(rx_en_dac), .I1(\rx_d[0] ), .O(data_to_dac)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7897.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7898 (.I0(\tx_dac_fsm_inst/sym_pos[0] ), .I1(\tx_dac_fsm_inst/sym_pos[1] ), 
            .O(\~tx_dac_fsm_inst/n431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__7898.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__7899 (.I0(\tx_dac_fsm_inst/sym_pos[0] ), .I1(\tx_dac_fsm_inst/sym_pos[1] ), 
            .I2(\tx_dac_fsm_inst/sym_pos[2] ), .O(\~tx_dac_fsm_inst/n436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__7899.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__7900 (.I0(\tx_dac_fsm_inst/sym_pos[0] ), .I1(\tx_dac_fsm_inst/sym_pos[1] ), 
            .I2(\tx_dac_fsm_inst/sym_pos[2] ), .I3(\tx_dac_fsm_inst/sym_pos[3] ), 
            .O(\~tx_dac_fsm_inst/n441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__7900.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__7901 (.I0(\tx_dac_fsm_inst/state_reg[2] ), .I1(\tx_dac_fsm_inst/zctr[1] ), 
            .I2(\tx_dac_fsm_inst/zctr[2] ), .I3(\tx_dac_fsm_inst/dac_config_reg[0] ), 
            .O(n4344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__7901.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__7902 (.I0(\tx_dac_fsm_inst/zctr[3] ), .I1(\tx_dac_fsm_inst/zctr[5] ), 
            .I2(\tx_dac_fsm_inst/zctr[4] ), .O(n4345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7902.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7903 (.I0(\tx_dac_fsm_inst/zctr[0] ), .I1(n4344), .I2(\tx_dac_fsm_inst/state_reg[0] ), 
            .I3(n4345), .O(n4346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__7903.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__7904 (.I0(n4335), .I1(\tx_dac_fsm_inst/state_reg[0] ), 
            .I2(n4346), .I3(\tx_dac_fsm_inst/state_reg[1] ), .O(n4347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__7904.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__7905 (.I0(n4342), .I1(n4332), .I2(n4347), .I3(\tx_dac_fsm_inst/state_reg[3] ), 
            .O(n3583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0 */ ;
    defparam LUT__7905.LUTMASK = 16'h88f0;
    EFX_LUT4 LUT__7906 (.I0(\tx_dac_fsm_inst/state_reg[0] ), .I1(\tx_dac_fsm_inst/state_reg[2] ), 
            .I2(n4331), .I3(\tx_dac_fsm_inst/state_reg[3] ), .O(n3584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__7906.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__7907 (.I0(n4333), .I1(\tx_dac_fsm_inst/state_reg[1] ), 
            .O(n3585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7907.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7908 (.I0(n4342), .I1(\tx_dac_fsm_inst/state_reg[3] ), 
            .I2(\tx_dac_fsm_inst/state_reg[0] ), .O(n3586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1818 */ ;
    defparam LUT__7908.LUTMASK = 16'h1818;
    EFX_LUT4 LUT__7909 (.I0(n115), .I1(n118), .O(\tx_dac_fsm_inst/n257 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7909.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7910 (.I0(n115), .I1(n3295), .O(\tx_dac_fsm_inst/n256 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7910.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7911 (.I0(n115), .I1(n3288), .O(\tx_dac_fsm_inst/n255 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7911.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7912 (.I0(n115), .I1(n3284), .O(\tx_dac_fsm_inst/n254 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7912.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7913 (.I0(n115), .I1(n3282), .O(\tx_dac_fsm_inst/n253 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7913.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7914 (.I0(n113), .I1(n121), .O(\tx_dac_fsm_inst/n283 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7914.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7915 (.I0(n113), .I1(n3276), .O(\tx_dac_fsm_inst/n282 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7915.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7916 (.I0(n113), .I1(n3273), .O(\tx_dac_fsm_inst/n281 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7916.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7917 (.I0(n113), .I1(n3269), .O(\tx_dac_fsm_inst/n280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7917.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7918 (.I0(n113), .I1(n3267), .O(\tx_dac_fsm_inst/n279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7918.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7919 (.I0(\reg_addr[4] ), .I1(n4343), .I2(n4240), .I3(\reg_addr[3] ), 
            .O(rx_en_fifo_length)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__7919.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__7920 (.I0(rx_en_fifo_length), .I1(\fifo_inst/wr_index[0] ), 
            .O(\fifo_inst/n153 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7920.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7921 (.I0(rx_en_fifo_length), .I1(n4319), .O(ceg_net146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7921.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7922 (.I0(rx_en_fifo_length), .I1(\fifo_inst/rd_index[0] ), 
            .O(\fifo_inst/n162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__7922.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__7923 (.I0(\fifo_inst/wr_index[0] ), .I1(\fifo_inst/rd_index[0] ), 
            .I2(\fifo_inst/wr_index[1] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__7923.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__7924 (.I0(\fifo_inst/wr_index[6] ), .I1(\fifo_inst/rd_index[6] ), 
            .I2(\fifo_inst/wr_index[7] ), .I3(\fifo_inst/rd_index[7] ), 
            .O(n4349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__7924.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__7925 (.I0(\fifo_inst/wr_index[2] ), .I1(\fifo_inst/rd_index[2] ), 
            .I2(\fifo_inst/wr_index[3] ), .I3(\fifo_inst/rd_index[3] ), 
            .O(n4350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__7925.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__7926 (.I0(\fifo_inst/wr_index[4] ), .I1(\fifo_inst/rd_index[4] ), 
            .I2(\fifo_inst/wr_index[5] ), .I3(\fifo_inst/rd_index[5] ), 
            .O(n4351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__7926.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__7927 (.I0(n4348), .I1(n4349), .I2(n4350), .I3(n4351), 
            .O(n4352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__7927.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__7928 (.I0(\fifo_inst/sync_rd[0] ), .I1(\fifo_inst/sync_rd[1] ), 
            .O(n4353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__7928.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__7929 (.I0(n4319), .I1(n4352), .I2(n4353), .I3(rx_en_fifo_length), 
            .O(ceg_net164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__7929.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__7930 (.I0(rx_en_fifo_length), .I1(\rx_d[0] ), .O(\data_to_fifo_length[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7930.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7931 (.I0(n4241), .I1(n4243), .O(tx_en_fifo)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__7931.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__7932 (.I0(\i14/fifo_inst/buff[20][0] ), .I1(\i14/fifo_inst/buff[22][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__7932.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__7933 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[1] ), 
            .I2(\fifo_inst/rd_index[2] ), .O(n4355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__7933.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__7934 (.I0(\i14/fifo_inst/buff[23][0] ), .I1(\i14/fifo_inst/buff[21][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7934.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7935 (.I0(n4354), .I1(n4356), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__7935.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__7936 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[1] ), 
            .I2(\fifo_inst/rd_index[3] ), .I3(\fifo_inst/rd_index[2] ), 
            .O(n4358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf78f */ ;
    defparam LUT__7936.LUTMASK = 16'hf78f;
    EFX_LUT4 LUT__7937 (.I0(\i14/fifo_inst/buff[24][0] ), .I1(\i14/fifo_inst/buff[26][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__7937.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__7938 (.I0(\i14/fifo_inst/buff[27][0] ), .I1(\i14/fifo_inst/buff[25][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7938.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7939 (.I0(n4358), .I1(n4359), .I2(n4360), .O(n4361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__7939.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__7940 (.I0(\i14/fifo_inst/buff[28][0] ), .I1(\i14/fifo_inst/buff[30][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__7940.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__7941 (.I0(\i14/fifo_inst/buff[31][0] ), .I1(\i14/fifo_inst/buff[29][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7941.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7942 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[1] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[3] ), 
            .O(n4364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__7942.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__7943 (.I0(n4362), .I1(n4363), .I2(n4364), .O(n4365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7943.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7944 (.I0(\i14/fifo_inst/buff[19][0] ), .I1(\i14/fifo_inst/buff[17][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7944.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7945 (.I0(\i14/fifo_inst/buff[16][0] ), .I1(\i14/fifo_inst/buff[18][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7945.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7946 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[1] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[3] ), 
            .O(n4368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ff8 */ ;
    defparam LUT__7946.LUTMASK = 16'h7ff8;
    EFX_LUT4 LUT__7947 (.I0(n4367), .I1(n4366), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7947.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7948 (.I0(n4357), .I1(n4361), .I2(n4365), .I3(n4369), 
            .O(n4370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__7948.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__7949 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[1] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[3] ), 
            .O(n4371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__7949.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__7950 (.I0(n4371), .I1(\fifo_inst/rd_index[4] ), .I2(\fifo_inst/rd_index[5] ), 
            .O(n4372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__7950.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__7951 (.I0(n4371), .I1(\fifo_inst/rd_index[4] ), .O(n4373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__7951.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__7952 (.I0(\i14/fifo_inst/buff[4][0] ), .I1(\i14/fifo_inst/buff[6][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__7952.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__7953 (.I0(\i14/fifo_inst/buff[7][0] ), .I1(\i14/fifo_inst/buff[5][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7953.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7954 (.I0(n4374), .I1(n4375), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__7954.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__7955 (.I0(\i14/fifo_inst/buff[12][0] ), .I1(\i14/fifo_inst/buff[14][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__7955.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__7956 (.I0(\i14/fifo_inst/buff[15][0] ), .I1(\i14/fifo_inst/buff[13][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7956.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7957 (.I0(n4377), .I1(n4378), .I2(n4364), .O(n4379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7957.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7958 (.I0(\i14/fifo_inst/buff[0][0] ), .I1(\i14/fifo_inst/buff[2][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__7958.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__7959 (.I0(\i14/fifo_inst/buff[3][0] ), .I1(\i14/fifo_inst/buff[1][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7959.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7960 (.I0(n4368), .I1(n4380), .I2(n4381), .O(n4382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__7960.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__7961 (.I0(\i14/fifo_inst/buff[8][0] ), .I1(\i14/fifo_inst/buff[10][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7961.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7962 (.I0(\i14/fifo_inst/buff[11][0] ), .I1(\i14/fifo_inst/buff[9][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7962.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7963 (.I0(n4384), .I1(n4383), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__7963.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__7964 (.I0(n4376), .I1(n4379), .I2(n4382), .I3(n4385), 
            .O(n4386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__7964.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__7965 (.I0(n4386), .I1(n4370), .I2(n4372), .I3(n4373), 
            .O(n4387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__7965.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__7966 (.I0(\i14/fifo_inst/buff[56][0] ), .I1(\i14/fifo_inst/buff[58][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7966.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7967 (.I0(\i14/fifo_inst/buff[59][0] ), .I1(\i14/fifo_inst/buff[57][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7967.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7968 (.I0(n4389), .I1(n4388), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__7968.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__7969 (.I0(\i14/fifo_inst/buff[52][0] ), .I1(\i14/fifo_inst/buff[54][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__7969.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__7970 (.I0(\i14/fifo_inst/buff[55][0] ), .I1(\i14/fifo_inst/buff[53][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7970.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7971 (.I0(n4391), .I1(n4392), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__7971.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__7972 (.I0(\i14/fifo_inst/buff[48][0] ), .I1(\i14/fifo_inst/buff[50][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__7972.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__7973 (.I0(\i14/fifo_inst/buff[51][0] ), .I1(\i14/fifo_inst/buff[49][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7973.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7974 (.I0(n4368), .I1(n4394), .I2(n4395), .O(n4396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__7974.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__7975 (.I0(\i14/fifo_inst/buff[60][0] ), .I1(\i14/fifo_inst/buff[62][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__7975.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__7976 (.I0(\i14/fifo_inst/buff[63][0] ), .I1(\i14/fifo_inst/buff[61][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7976.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7977 (.I0(n4397), .I1(n4398), .I2(n4364), .O(n4399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7977.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7978 (.I0(n4390), .I1(n4393), .I2(n4396), .I3(n4399), 
            .O(n4400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__7978.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__7979 (.I0(\i14/fifo_inst/buff[32][0] ), .I1(\i14/fifo_inst/buff[34][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__7979.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__7980 (.I0(\i14/fifo_inst/buff[35][0] ), .I1(\i14/fifo_inst/buff[33][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7980.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7981 (.I0(n4368), .I1(n4401), .I2(n4402), .O(n4403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__7981.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__7982 (.I0(\i14/fifo_inst/buff[44][0] ), .I1(\i14/fifo_inst/buff[46][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__7982.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__7983 (.I0(\i14/fifo_inst/buff[47][0] ), .I1(\i14/fifo_inst/buff[45][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7983.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7984 (.I0(n4404), .I1(n4405), .I2(n4364), .O(n4406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__7984.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__7985 (.I0(\i14/fifo_inst/buff[40][0] ), .I1(\i14/fifo_inst/buff[42][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7985.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7986 (.I0(\i14/fifo_inst/buff[43][0] ), .I1(\i14/fifo_inst/buff[41][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7986.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7987 (.I0(n4408), .I1(n4407), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__7987.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__7988 (.I0(\i14/fifo_inst/buff[36][0] ), .I1(\i14/fifo_inst/buff[38][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__7988.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__7989 (.I0(\i14/fifo_inst/buff[39][0] ), .I1(\i14/fifo_inst/buff[37][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7989.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7990 (.I0(n4410), .I1(n4411), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__7990.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__7991 (.I0(n4403), .I1(n4406), .I2(n4409), .I3(n4412), 
            .O(n4413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__7991.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__7992 (.I0(n4413), .I1(n4400), .I2(n4372), .I3(n4387), 
            .O(n4414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3f50 */ ;
    defparam LUT__7992.LUTMASK = 16'h3f50;
    EFX_LUT4 LUT__7993 (.I0(n4371), .I1(\fifo_inst/rd_index[4] ), .I2(\fifo_inst/rd_index[5] ), 
            .O(n4415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__7993.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__7994 (.I0(n4415), .I1(\fifo_inst/rd_index[6] ), .O(n4416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__7994.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__7995 (.I0(\i14/fifo_inst/buff[68][0] ), .I1(\i14/fifo_inst/buff[70][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__7995.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__7996 (.I0(\i14/fifo_inst/buff[71][0] ), .I1(\i14/fifo_inst/buff[69][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__7996.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__7997 (.I0(n4417), .I1(n4418), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__7997.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__7998 (.I0(\i14/fifo_inst/buff[76][0] ), .I1(\i14/fifo_inst/buff[78][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7998.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__7999 (.I0(\i14/fifo_inst/buff[79][0] ), .I1(\i14/fifo_inst/buff[77][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__7999.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8000 (.I0(n4421), .I1(n4420), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4364), .O(n4422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8000.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8001 (.I0(\i14/fifo_inst/buff[75][0] ), .I1(\i14/fifo_inst/buff[73][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8001.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8002 (.I0(\i14/fifo_inst/buff[72][0] ), .I1(\i14/fifo_inst/buff[74][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8002.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8003 (.I0(n4424), .I1(n4423), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8003.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8004 (.I0(\i14/fifo_inst/buff[64][0] ), .I1(\i14/fifo_inst/buff[66][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8004.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8005 (.I0(\i14/fifo_inst/buff[67][0] ), .I1(\i14/fifo_inst/buff[65][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8005.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8006 (.I0(n4427), .I1(n4426), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8006.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8007 (.I0(n4419), .I1(n4422), .I2(n4425), .I3(n4428), 
            .O(n4429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8007.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8008 (.I0(\i14/fifo_inst/buff[100][0] ), .I1(\i14/fifo_inst/buff[101][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haffc */ ;
    defparam LUT__8008.LUTMASK = 16'haffc;
    EFX_LUT4 LUT__8009 (.I0(\i14/fifo_inst/buff[102][0] ), .I1(\i14/fifo_inst/buff[103][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfacf */ ;
    defparam LUT__8009.LUTMASK = 16'hfacf;
    EFX_LUT4 LUT__8010 (.I0(\fifo_inst/rd_index[3] ), .I1(n4355), .I2(n4430), 
            .I3(n4431), .O(n4432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__8010.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__8011 (.I0(\i14/fifo_inst/buff[96][0] ), .I1(\i14/fifo_inst/buff[98][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8011.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8012 (.I0(\i14/fifo_inst/buff[99][0] ), .I1(\i14/fifo_inst/buff[97][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8012.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8013 (.I0(n4434), .I1(n4433), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8013.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8014 (.I0(\i14/fifo_inst/buff[107][0] ), .I1(\i14/fifo_inst/buff[105][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8014.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8015 (.I0(\i14/fifo_inst/buff[104][0] ), .I1(\i14/fifo_inst/buff[106][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8015.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8016 (.I0(n4358), .I1(n4436), .I2(n4437), .O(n4438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8016.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8017 (.I0(\i14/fifo_inst/buff[108][0] ), .I1(\i14/fifo_inst/buff[110][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8017.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8018 (.I0(\i14/fifo_inst/buff[111][0] ), .I1(\i14/fifo_inst/buff[109][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8018.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8019 (.I0(n4439), .I1(n4440), .I2(n4364), .O(n4441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8019.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8020 (.I0(n4432), .I1(n4435), .I2(n4438), .I3(n4441), 
            .O(n4442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8020.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8021 (.I0(n4442), .I1(n4429), .I2(n4373), .I3(n4372), 
            .O(n4443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8021.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8022 (.I0(\i14/fifo_inst/buff[112][0] ), .I1(\i14/fifo_inst/buff[114][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8022.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8023 (.I0(\i14/fifo_inst/buff[115][0] ), .I1(\i14/fifo_inst/buff[113][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8023.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8024 (.I0(n4368), .I1(n4444), .I2(n4445), .O(n4446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8024.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8025 (.I0(\i14/fifo_inst/buff[120][0] ), .I1(\i14/fifo_inst/buff[122][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8025.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8026 (.I0(\i14/fifo_inst/buff[123][0] ), .I1(\i14/fifo_inst/buff[121][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8026.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8027 (.I0(n4448), .I1(n4447), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8027.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8028 (.I0(\i14/fifo_inst/buff[116][0] ), .I1(\i14/fifo_inst/buff[118][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8028.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8029 (.I0(\i14/fifo_inst/buff[119][0] ), .I1(\i14/fifo_inst/buff[117][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8029.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8030 (.I0(n4450), .I1(n4451), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8030.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8031 (.I0(\i14/fifo_inst/buff[124][0] ), .I1(\i14/fifo_inst/buff[126][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8031.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8032 (.I0(\i14/fifo_inst/buff[127][0] ), .I1(\i14/fifo_inst/buff[125][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8032.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8033 (.I0(n4453), .I1(n4454), .I2(n4364), .O(n4455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8033.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8034 (.I0(n4446), .I1(n4449), .I2(n4452), .I3(n4455), 
            .O(n4456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8034.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8035 (.I0(\i14/fifo_inst/buff[84][0] ), .I1(\i14/fifo_inst/buff[86][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8035.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8036 (.I0(\i14/fifo_inst/buff[87][0] ), .I1(\i14/fifo_inst/buff[85][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8036.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8037 (.I0(n4457), .I1(n4458), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8037.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8038 (.I0(\i14/fifo_inst/buff[88][0] ), .I1(\i14/fifo_inst/buff[90][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8038.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8039 (.I0(\i14/fifo_inst/buff[91][0] ), .I1(\i14/fifo_inst/buff[89][0] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8039.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8040 (.I0(n4358), .I1(n4460), .I2(n4461), .O(n4462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8040.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8041 (.I0(\i14/fifo_inst/buff[92][0] ), .I1(\i14/fifo_inst/buff[94][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8041.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8042 (.I0(\i14/fifo_inst/buff[95][0] ), .I1(\i14/fifo_inst/buff[93][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8042.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8043 (.I0(n4464), .I1(n4463), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4364), .O(n4465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8043.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8044 (.I0(\i14/fifo_inst/buff[83][0] ), .I1(\i14/fifo_inst/buff[81][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8044.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8045 (.I0(\i14/fifo_inst/buff[80][0] ), .I1(\i14/fifo_inst/buff[82][0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8045.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8046 (.I0(n4467), .I1(n4466), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8046.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8047 (.I0(n4459), .I1(n4462), .I2(n4465), .I3(n4468), 
            .O(n4469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8047.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8048 (.I0(n4469), .I1(n4456), .I2(n4372), .I3(n4373), 
            .O(n4470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8048.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8049 (.I0(n4352), .I1(ceg_net146), .O(n4471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8049.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8050 (.I0(n4443), .I1(n4470), .I2(n4416), .I3(n4471), 
            .O(n4472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8050.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8051 (.I0(n4319), .I1(n4416), .O(n4473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8051.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8052 (.I0(rx_en_fifo), .I1(n4319), .I2(\rx_d[0] ), .O(n4474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__8052.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__8053 (.I0(n4472), .I1(n4474), .I2(n4414), .I3(n4473), 
            .O(\fifo_inst/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__8053.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__8054 (.I0(n4353), .I1(rx_en_fifo_length), .I2(n4352), 
            .I3(n4319), .O(ceg_net418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f11 */ ;
    defparam LUT__8054.LUTMASK = 16'h0f11;
    EFX_LUT4 LUT__8055 (.I0(rx_en_fifo_length), .I1(n124), .O(\fifo_inst/n152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8055.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8056 (.I0(rx_en_fifo_length), .I1(n3260), .O(\fifo_inst/n151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8056.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8057 (.I0(rx_en_fifo_length), .I1(n3237), .O(\fifo_inst/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8057.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8058 (.I0(rx_en_fifo_length), .I1(n3234), .O(\fifo_inst/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8058.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8059 (.I0(rx_en_fifo_length), .I1(n3231), .O(\fifo_inst/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8059.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8060 (.I0(rx_en_fifo_length), .I1(n3228), .O(\fifo_inst/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8060.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8061 (.I0(rx_en_fifo_length), .I1(n3226), .O(\fifo_inst/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8061.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8062 (.I0(rx_en_fifo_length), .I1(\fifo_inst/rd_index[0] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(\fifo_inst/n161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__8062.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__8063 (.I0(rx_en_fifo_length), .I1(n4355), .O(\fifo_inst/n160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8063.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8064 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[1] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\fifo_inst/rd_index[3] ), 
            .O(n4475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h807f */ ;
    defparam LUT__8064.LUTMASK = 16'h807f;
    EFX_LUT4 LUT__8065 (.I0(rx_en_fifo_length), .I1(n4475), .O(\fifo_inst/n159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8065.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8066 (.I0(rx_en_fifo_length), .I1(n4373), .O(\fifo_inst/n158 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8066.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8067 (.I0(rx_en_fifo_length), .I1(n4372), .O(\fifo_inst/n157 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8067.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8068 (.I0(rx_en_fifo_length), .I1(n4416), .O(\fifo_inst/n156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8068.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8069 (.I0(n4415), .I1(\fifo_inst/rd_index[6] ), .I2(rx_en_fifo_length), 
            .I3(\fifo_inst/rd_index[7] ), .O(\fifo_inst/n155 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__8069.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__8070 (.I0(rx_en_fifo_length), .I1(\rx_d[1] ), .O(\data_to_fifo_length[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8070.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8071 (.I0(rx_en_fifo_length), .I1(\rx_d[2] ), .O(\data_to_fifo_length[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8071.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8072 (.I0(rx_en_fifo_length), .I1(\rx_d[3] ), .O(\data_to_fifo_length[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8072.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8073 (.I0(rx_en_fifo_length), .I1(\rx_d[4] ), .O(\data_to_fifo_length[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8073.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8074 (.I0(rx_en_fifo_length), .I1(\rx_d[5] ), .O(\data_to_fifo_length[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8074.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8075 (.I0(rx_en_fifo_length), .I1(\rx_d[6] ), .O(\data_to_fifo_length[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8075.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8076 (.I0(rx_en_fifo_length), .I1(\rx_d[7] ), .O(\data_to_fifo_length[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8076.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8077 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[2] ), 
            .I2(\fifo_inst/wr_index[3] ), .I3(\fifo_inst/wr_index[4] ), 
            .O(n4476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8077.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8078 (.I0(n4324), .I1(n4476), .O(\i14/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8078.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8079 (.I0(rx_en_fifo), .I1(\rx_d[4] ), .O(\data_to_fifo[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8079.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8080 (.I0(n4321), .I1(n4476), .O(\i14/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8080.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8081 (.I0(rx_en_fifo), .I1(\rx_d[5] ), .O(\data_to_fifo[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8081.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8082 (.I0(rx_en_fifo), .I1(\rx_d[3] ), .O(\data_to_fifo[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8082.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8083 (.I0(rx_en_fifo), .I1(n4319), .I2(\rx_d[1] ), .O(n4477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__8083.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__8084 (.I0(\i14/fifo_inst/buff[63][1] ), .I1(\i14/fifo_inst/buff[61][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8084.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8085 (.I0(\i14/fifo_inst/buff[60][1] ), .I1(\i14/fifo_inst/buff[62][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8085.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8086 (.I0(n4478), .I1(n4479), .I2(n4364), .O(n4480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8086.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8087 (.I0(\i14/fifo_inst/buff[56][1] ), .I1(\i14/fifo_inst/buff[57][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haffc */ ;
    defparam LUT__8087.LUTMASK = 16'haffc;
    EFX_LUT4 LUT__8088 (.I0(\i14/fifo_inst/buff[58][1] ), .I1(\i14/fifo_inst/buff[59][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfacf */ ;
    defparam LUT__8088.LUTMASK = 16'hfacf;
    EFX_LUT4 LUT__8089 (.I0(n4358), .I1(n4481), .I2(n4482), .O(n4483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__8089.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__8090 (.I0(\i14/fifo_inst/buff[48][1] ), .I1(\i14/fifo_inst/buff[50][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8090.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8091 (.I0(\i14/fifo_inst/buff[51][1] ), .I1(\i14/fifo_inst/buff[49][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8091.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8092 (.I0(n4485), .I1(n4484), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8092.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8093 (.I0(\i14/fifo_inst/buff[55][1] ), .I1(\i14/fifo_inst/buff[53][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8093.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8094 (.I0(\i14/fifo_inst/buff[52][1] ), .I1(\i14/fifo_inst/buff[54][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8094.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8095 (.I0(n4487), .I1(n4488), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8095.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8096 (.I0(n4480), .I1(n4483), .I2(n4486), .I3(n4489), 
            .O(n4490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8096.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8097 (.I0(\i14/fifo_inst/buff[28][1] ), .I1(\i14/fifo_inst/buff[30][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8097.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8098 (.I0(\i14/fifo_inst/buff[31][1] ), .I1(\i14/fifo_inst/buff[29][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8098.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8099 (.I0(n4492), .I1(n4491), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4364), .O(n4493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8099.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8100 (.I0(\i14/fifo_inst/buff[20][1] ), .I1(\i14/fifo_inst/buff[22][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8100.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8101 (.I0(\i14/fifo_inst/buff[23][1] ), .I1(\i14/fifo_inst/buff[21][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8101.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8102 (.I0(n4494), .I1(n4495), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8102.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8103 (.I0(\i14/fifo_inst/buff[24][1] ), .I1(\i14/fifo_inst/buff[26][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8103.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8104 (.I0(\i14/fifo_inst/buff[27][1] ), .I1(\i14/fifo_inst/buff[25][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8104.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8105 (.I0(n4358), .I1(n4497), .I2(n4498), .O(n4499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8105.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8106 (.I0(\i14/fifo_inst/buff[16][1] ), .I1(\i14/fifo_inst/buff[17][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haffc */ ;
    defparam LUT__8106.LUTMASK = 16'haffc;
    EFX_LUT4 LUT__8107 (.I0(\i14/fifo_inst/buff[18][1] ), .I1(\i14/fifo_inst/buff[19][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfacf */ ;
    defparam LUT__8107.LUTMASK = 16'hfacf;
    EFX_LUT4 LUT__8108 (.I0(n4368), .I1(n4500), .I2(n4501), .O(n4502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__8108.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__8109 (.I0(n4493), .I1(n4496), .I2(n4499), .I3(n4502), 
            .O(n4503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8109.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8110 (.I0(n4503), .I1(n4490), .I2(n4372), .I3(n4373), 
            .O(n4504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8110.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8111 (.I0(\i14/fifo_inst/buff[32][1] ), .I1(\i14/fifo_inst/buff[34][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8111.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8112 (.I0(\i14/fifo_inst/buff[35][1] ), .I1(\i14/fifo_inst/buff[33][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8112.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8113 (.I0(n4506), .I1(n4505), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8113.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8114 (.I0(\i14/fifo_inst/buff[36][1] ), .I1(\i14/fifo_inst/buff[38][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8114.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8115 (.I0(\i14/fifo_inst/buff[39][1] ), .I1(\i14/fifo_inst/buff[37][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8115.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8116 (.I0(n4508), .I1(n4509), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8116.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8117 (.I0(\i14/fifo_inst/buff[40][1] ), .I1(\i14/fifo_inst/buff[42][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8117.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8118 (.I0(\i14/fifo_inst/buff[43][1] ), .I1(\i14/fifo_inst/buff[41][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8118.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8119 (.I0(n4512), .I1(n4511), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8119.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8120 (.I0(\i14/fifo_inst/buff[44][1] ), .I1(\i14/fifo_inst/buff[46][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8120.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8121 (.I0(\i14/fifo_inst/buff[47][1] ), .I1(\i14/fifo_inst/buff[45][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8121.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8122 (.I0(n4514), .I1(n4515), .I2(n4364), .O(n4516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8122.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8123 (.I0(n4507), .I1(n4510), .I2(n4513), .I3(n4516), 
            .O(n4517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8123.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8124 (.I0(\i14/fifo_inst/buff[4][1] ), .I1(\i14/fifo_inst/buff[6][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8124.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8125 (.I0(\i14/fifo_inst/buff[7][1] ), .I1(\i14/fifo_inst/buff[5][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8125.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8126 (.I0(n4518), .I1(n4519), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8126.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8127 (.I0(\i14/fifo_inst/buff[8][1] ), .I1(\i14/fifo_inst/buff[10][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8127.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8128 (.I0(\i14/fifo_inst/buff[11][1] ), .I1(\i14/fifo_inst/buff[9][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8128.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8129 (.I0(n4522), .I1(n4521), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8129.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8130 (.I0(\i14/fifo_inst/buff[12][1] ), .I1(\i14/fifo_inst/buff[14][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8130.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8131 (.I0(\i14/fifo_inst/buff[15][1] ), .I1(\i14/fifo_inst/buff[13][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8131.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8132 (.I0(n4524), .I1(n4525), .I2(n4364), .O(n4526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8132.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8133 (.I0(\i14/fifo_inst/buff[3][1] ), .I1(\i14/fifo_inst/buff[1][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8133.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8134 (.I0(\i14/fifo_inst/buff[0][1] ), .I1(\i14/fifo_inst/buff[2][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8134.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8135 (.I0(n4528), .I1(n4527), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8135.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8136 (.I0(n4520), .I1(n4523), .I2(n4526), .I3(n4529), 
            .O(n4530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8136.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8137 (.I0(n4530), .I1(n4517), .I2(n4373), .I3(n4372), 
            .O(n4531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8137.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8138 (.I0(n4504), .I1(n4531), .I2(n4477), .I3(n4416), 
            .O(n4532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8138.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8139 (.I0(\i14/fifo_inst/buff[84][1] ), .I1(\i14/fifo_inst/buff[86][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8139.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8140 (.I0(\i14/fifo_inst/buff[87][1] ), .I1(\i14/fifo_inst/buff[85][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8140.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8141 (.I0(n4533), .I1(n4534), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8141.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8142 (.I0(\i14/fifo_inst/buff[92][1] ), .I1(\i14/fifo_inst/buff[94][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8142.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8143 (.I0(\i14/fifo_inst/buff[95][1] ), .I1(\i14/fifo_inst/buff[93][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8143.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8144 (.I0(n4536), .I1(n4537), .I2(n4364), .O(n4538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8144.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8145 (.I0(\i14/fifo_inst/buff[88][1] ), .I1(\i14/fifo_inst/buff[90][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8145.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8146 (.I0(\i14/fifo_inst/buff[91][1] ), .I1(\i14/fifo_inst/buff[89][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8146.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8147 (.I0(n4358), .I1(n4539), .I2(n4540), .O(n4541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8147.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8148 (.I0(\i14/fifo_inst/buff[80][1] ), .I1(\i14/fifo_inst/buff[82][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8148.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8149 (.I0(\i14/fifo_inst/buff[83][1] ), .I1(\i14/fifo_inst/buff[81][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8149.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8150 (.I0(n4543), .I1(n4542), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8150.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8151 (.I0(n4535), .I1(n4538), .I2(n4541), .I3(n4544), 
            .O(n4545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8151.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8152 (.I0(\i14/fifo_inst/buff[124][1] ), .I1(\i14/fifo_inst/buff[126][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8152.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8153 (.I0(\i14/fifo_inst/buff[127][1] ), .I1(\i14/fifo_inst/buff[125][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8153.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8154 (.I0(n4547), .I1(n4546), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4364), .O(n4548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8154.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8155 (.I0(\i14/fifo_inst/buff[116][1] ), .I1(\i14/fifo_inst/buff[118][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8155.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8156 (.I0(\i14/fifo_inst/buff[119][1] ), .I1(\i14/fifo_inst/buff[117][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8156.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8157 (.I0(n4549), .I1(n4550), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8157.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8158 (.I0(\i14/fifo_inst/buff[120][1] ), .I1(\i14/fifo_inst/buff[122][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8158.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8159 (.I0(\i14/fifo_inst/buff[123][1] ), .I1(\i14/fifo_inst/buff[121][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8159.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8160 (.I0(n4553), .I1(n4552), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8160.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8161 (.I0(\i14/fifo_inst/buff[112][1] ), .I1(\i14/fifo_inst/buff[114][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8161.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8162 (.I0(\i14/fifo_inst/buff[115][1] ), .I1(\i14/fifo_inst/buff[113][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8162.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8163 (.I0(n4556), .I1(n4555), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8163.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8164 (.I0(n4548), .I1(n4551), .I2(n4554), .I3(n4557), 
            .O(n4558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8164.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8165 (.I0(n4558), .I1(n4545), .I2(n4372), .I3(n4373), 
            .O(n4559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8165.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8166 (.I0(\i14/fifo_inst/buff[68][1] ), .I1(\i14/fifo_inst/buff[70][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8166.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8167 (.I0(\i14/fifo_inst/buff[71][1] ), .I1(\i14/fifo_inst/buff[69][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8167.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8168 (.I0(n4560), .I1(n4561), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8168.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8169 (.I0(\i14/fifo_inst/buff[72][1] ), .I1(\i14/fifo_inst/buff[74][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8169.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8170 (.I0(\i14/fifo_inst/buff[75][1] ), .I1(\i14/fifo_inst/buff[73][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8170.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8171 (.I0(n4564), .I1(n4563), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8171.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8172 (.I0(\i14/fifo_inst/buff[76][1] ), .I1(\i14/fifo_inst/buff[78][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8172.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8173 (.I0(\i14/fifo_inst/buff[79][1] ), .I1(\i14/fifo_inst/buff[77][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8173.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8174 (.I0(n4566), .I1(n4567), .I2(n4364), .O(n4568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8174.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8175 (.I0(\i14/fifo_inst/buff[67][1] ), .I1(\i14/fifo_inst/buff[65][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8175.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8176 (.I0(\i14/fifo_inst/buff[64][1] ), .I1(\i14/fifo_inst/buff[66][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8176.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8177 (.I0(n4570), .I1(n4569), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8177.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8178 (.I0(n4562), .I1(n4565), .I2(n4568), .I3(n4571), 
            .O(n4572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8178.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8179 (.I0(\i14/fifo_inst/buff[96][1] ), .I1(\i14/fifo_inst/buff[98][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8179.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8180 (.I0(\i14/fifo_inst/buff[99][1] ), .I1(\i14/fifo_inst/buff[97][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8180.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8181 (.I0(n4368), .I1(n4573), .I2(n4574), .O(n4575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8181.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8182 (.I0(\i14/fifo_inst/buff[104][1] ), .I1(\i14/fifo_inst/buff[106][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8182.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8183 (.I0(\i14/fifo_inst/buff[107][1] ), .I1(\i14/fifo_inst/buff[105][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8183.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8184 (.I0(n4577), .I1(n4576), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8184.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8185 (.I0(\i14/fifo_inst/buff[108][1] ), .I1(\i14/fifo_inst/buff[110][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8185.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8186 (.I0(\i14/fifo_inst/buff[111][1] ), .I1(\i14/fifo_inst/buff[109][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8186.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8187 (.I0(n4580), .I1(n4579), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4364), .O(n4581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8187.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8188 (.I0(\i14/fifo_inst/buff[100][1] ), .I1(\i14/fifo_inst/buff[102][1] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8188.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8189 (.I0(\i14/fifo_inst/buff[103][1] ), .I1(\i14/fifo_inst/buff[101][1] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8189.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8190 (.I0(n4582), .I1(n4583), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8190.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8191 (.I0(n4575), .I1(n4578), .I2(n4581), .I3(n4584), 
            .O(n4585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8191.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8192 (.I0(n4585), .I1(n4572), .I2(n4373), .I3(n4372), 
            .O(n4586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8192.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8193 (.I0(n4477), .I1(n4559), .I2(n4586), .I3(n4416), 
            .O(n4587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8193.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8194 (.I0(n4471), .I1(n4477), .I2(n4532), .I3(n4587), 
            .O(\fifo_inst/n143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__8194.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__8195 (.I0(rx_en_fifo), .I1(n4319), .I2(\rx_d[2] ), .O(n4588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__8195.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__8196 (.I0(\i14/fifo_inst/buff[11][2] ), .I1(\i14/fifo_inst/buff[9][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8196.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8197 (.I0(\i14/fifo_inst/buff[8][2] ), .I1(\i14/fifo_inst/buff[10][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8197.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8198 (.I0(n4358), .I1(n4589), .I2(n4590), .O(n4591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8198.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8199 (.I0(\i14/fifo_inst/buff[4][2] ), .I1(\i14/fifo_inst/buff[6][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8199.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8200 (.I0(\i14/fifo_inst/buff[7][2] ), .I1(\i14/fifo_inst/buff[5][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8200.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8201 (.I0(n4592), .I1(n4593), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8201.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8202 (.I0(\i14/fifo_inst/buff[12][2] ), .I1(\i14/fifo_inst/buff[14][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8202.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8203 (.I0(\i14/fifo_inst/buff[15][2] ), .I1(\i14/fifo_inst/buff[13][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8203.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8204 (.I0(n4596), .I1(n4595), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4364), .O(n4597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8204.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8205 (.I0(\i14/fifo_inst/buff[3][2] ), .I1(\i14/fifo_inst/buff[1][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8205.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8206 (.I0(\i14/fifo_inst/buff[0][2] ), .I1(\i14/fifo_inst/buff[2][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8206.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8207 (.I0(n4599), .I1(n4598), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8207.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8208 (.I0(n4591), .I1(n4594), .I2(n4597), .I3(n4600), 
            .O(n4601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8208.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8209 (.I0(\i14/fifo_inst/buff[36][2] ), .I1(\i14/fifo_inst/buff[38][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8209.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8210 (.I0(\i14/fifo_inst/buff[39][2] ), .I1(\i14/fifo_inst/buff[37][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8210.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8211 (.I0(n4602), .I1(n4603), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8211.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8212 (.I0(\i14/fifo_inst/buff[40][2] ), .I1(\i14/fifo_inst/buff[42][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8212.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8213 (.I0(\i14/fifo_inst/buff[43][2] ), .I1(\i14/fifo_inst/buff[41][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8213.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8214 (.I0(n4606), .I1(n4605), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8214.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8215 (.I0(\i14/fifo_inst/buff[32][2] ), .I1(\i14/fifo_inst/buff[34][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8215.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8216 (.I0(\i14/fifo_inst/buff[35][2] ), .I1(\i14/fifo_inst/buff[33][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8216.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8217 (.I0(n4368), .I1(n4608), .I2(n4609), .O(n4610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8217.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8218 (.I0(\i14/fifo_inst/buff[44][2] ), .I1(\i14/fifo_inst/buff[46][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8218.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8219 (.I0(\i14/fifo_inst/buff[47][2] ), .I1(\i14/fifo_inst/buff[45][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8219.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8220 (.I0(n4611), .I1(n4612), .I2(n4364), .O(n4613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8220.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8221 (.I0(n4604), .I1(n4607), .I2(n4610), .I3(n4613), 
            .O(n4614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8221.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8222 (.I0(n4614), .I1(n4601), .I2(n4373), .I3(n4372), 
            .O(n4615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8222.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8223 (.I0(\i14/fifo_inst/buff[60][2] ), .I1(\i14/fifo_inst/buff[62][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8223.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8224 (.I0(\i14/fifo_inst/buff[63][2] ), .I1(\i14/fifo_inst/buff[61][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8224.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8225 (.I0(n4616), .I1(n4617), .I2(n4364), .O(n4618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8225.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8226 (.I0(\i14/fifo_inst/buff[48][2] ), .I1(\i14/fifo_inst/buff[50][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4619)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8226.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8227 (.I0(\i14/fifo_inst/buff[51][2] ), .I1(\i14/fifo_inst/buff[49][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8227.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8228 (.I0(n4368), .I1(n4619), .I2(n4620), .O(n4621)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8228.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8229 (.I0(\i14/fifo_inst/buff[52][2] ), .I1(\i14/fifo_inst/buff[54][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8229.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8230 (.I0(\i14/fifo_inst/buff[55][2] ), .I1(\i14/fifo_inst/buff[53][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8230.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8231 (.I0(n4622), .I1(n4623), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8231.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8232 (.I0(\i14/fifo_inst/buff[56][2] ), .I1(\i14/fifo_inst/buff[58][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8232.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8233 (.I0(\i14/fifo_inst/buff[59][2] ), .I1(\i14/fifo_inst/buff[57][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8233.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8234 (.I0(n4626), .I1(n4625), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8234.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8235 (.I0(n4618), .I1(n4621), .I2(n4624), .I3(n4627), 
            .O(n4628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8235.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8236 (.I0(\i14/fifo_inst/buff[20][2] ), .I1(\i14/fifo_inst/buff[22][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8236.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8237 (.I0(\i14/fifo_inst/buff[23][2] ), .I1(\i14/fifo_inst/buff[21][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8237.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8238 (.I0(n4629), .I1(n4630), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8238.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8239 (.I0(\i14/fifo_inst/buff[24][2] ), .I1(\i14/fifo_inst/buff[26][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8239.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8240 (.I0(\i14/fifo_inst/buff[27][2] ), .I1(\i14/fifo_inst/buff[25][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8240.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8241 (.I0(n4358), .I1(n4632), .I2(n4633), .O(n4634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8241.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8242 (.I0(\i14/fifo_inst/buff[28][2] ), .I1(\i14/fifo_inst/buff[30][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8242.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8243 (.I0(\i14/fifo_inst/buff[31][2] ), .I1(\i14/fifo_inst/buff[29][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8243.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8244 (.I0(n4636), .I1(n4635), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4364), .O(n4637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8244.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8245 (.I0(\i14/fifo_inst/buff[16][2] ), .I1(\i14/fifo_inst/buff[18][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8245.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8246 (.I0(\i14/fifo_inst/buff[19][2] ), .I1(\i14/fifo_inst/buff[17][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8246.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8247 (.I0(n4639), .I1(n4638), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4640)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8247.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8248 (.I0(n4631), .I1(n4634), .I2(n4637), .I3(n4640), 
            .O(n4641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8248.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8249 (.I0(n4641), .I1(n4628), .I2(n4372), .I3(n4373), 
            .O(n4642)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8249.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8250 (.I0(n4615), .I1(n4588), .I2(n4642), .I3(n4416), 
            .O(n4643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8250.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8251 (.I0(\i14/fifo_inst/buff[76][2] ), .I1(\i14/fifo_inst/buff[78][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8251.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8252 (.I0(\i14/fifo_inst/buff[79][2] ), .I1(\i14/fifo_inst/buff[77][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8252.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8253 (.I0(n4645), .I1(n4644), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4364), .O(n4646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8253.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8254 (.I0(\i14/fifo_inst/buff[68][2] ), .I1(\i14/fifo_inst/buff[70][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8254.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8255 (.I0(\i14/fifo_inst/buff[71][2] ), .I1(\i14/fifo_inst/buff[69][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8255.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8256 (.I0(n4647), .I1(n4648), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8256.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8257 (.I0(\i14/fifo_inst/buff[75][2] ), .I1(\i14/fifo_inst/buff[73][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8257.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8258 (.I0(\i14/fifo_inst/buff[72][2] ), .I1(\i14/fifo_inst/buff[74][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8258.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8259 (.I0(n4651), .I1(n4650), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8259.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8260 (.I0(\i14/fifo_inst/buff[64][2] ), .I1(\i14/fifo_inst/buff[66][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8260.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8261 (.I0(\i14/fifo_inst/buff[67][2] ), .I1(\i14/fifo_inst/buff[65][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8261.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8262 (.I0(n4654), .I1(n4653), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8262.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8263 (.I0(n4646), .I1(n4649), .I2(n4652), .I3(n4655), 
            .O(n4656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8263.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8264 (.I0(\i14/fifo_inst/buff[108][2] ), .I1(\i14/fifo_inst/buff[110][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8264.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8265 (.I0(\i14/fifo_inst/buff[111][2] ), .I1(\i14/fifo_inst/buff[109][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8265.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8266 (.I0(n4658), .I1(n4657), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4364), .O(n4659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8266.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8267 (.I0(\i14/fifo_inst/buff[96][2] ), .I1(\i14/fifo_inst/buff[98][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8267.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8268 (.I0(\i14/fifo_inst/buff[99][2] ), .I1(\i14/fifo_inst/buff[97][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8268.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8269 (.I0(n4661), .I1(n4660), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8269.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8270 (.I0(\i14/fifo_inst/buff[100][2] ), .I1(\i14/fifo_inst/buff[102][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8270.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8271 (.I0(\i14/fifo_inst/buff[103][2] ), .I1(\i14/fifo_inst/buff[101][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8271.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8272 (.I0(n4663), .I1(n4664), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8272.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8273 (.I0(\i14/fifo_inst/buff[104][2] ), .I1(\i14/fifo_inst/buff[106][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8273.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8274 (.I0(\i14/fifo_inst/buff[107][2] ), .I1(\i14/fifo_inst/buff[105][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8274.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8275 (.I0(n4667), .I1(n4666), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8275.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8276 (.I0(n4659), .I1(n4662), .I2(n4665), .I3(n4668), 
            .O(n4669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8276.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8277 (.I0(n4669), .I1(n4656), .I2(n4373), .I3(n4372), 
            .O(n4670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8277.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8278 (.I0(\i14/fifo_inst/buff[80][2] ), .I1(\i14/fifo_inst/buff[82][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8278.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8279 (.I0(\i14/fifo_inst/buff[83][2] ), .I1(\i14/fifo_inst/buff[81][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8279.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8280 (.I0(n4368), .I1(n4671), .I2(n4672), .O(n4673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8280.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8281 (.I0(\i14/fifo_inst/buff[88][2] ), .I1(\i14/fifo_inst/buff[90][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8281.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8282 (.I0(\i14/fifo_inst/buff[91][2] ), .I1(\i14/fifo_inst/buff[89][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8282.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8283 (.I0(n4675), .I1(n4674), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8283.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8284 (.I0(\i14/fifo_inst/buff[92][2] ), .I1(\i14/fifo_inst/buff[94][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4677)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8284.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8285 (.I0(\i14/fifo_inst/buff[95][2] ), .I1(\i14/fifo_inst/buff[93][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8285.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8286 (.I0(n4678), .I1(n4677), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4364), .O(n4679)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8286.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8287 (.I0(\i14/fifo_inst/buff[84][2] ), .I1(\i14/fifo_inst/buff[86][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8287.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8288 (.I0(\i14/fifo_inst/buff[87][2] ), .I1(\i14/fifo_inst/buff[85][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4681)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8288.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8289 (.I0(n4680), .I1(n4681), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8289.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8290 (.I0(n4673), .I1(n4676), .I2(n4679), .I3(n4682), 
            .O(n4683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8290.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8291 (.I0(\i14/fifo_inst/buff[112][2] ), .I1(\i14/fifo_inst/buff[114][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8291.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8292 (.I0(\i14/fifo_inst/buff[115][2] ), .I1(\i14/fifo_inst/buff[113][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8292.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8293 (.I0(n4685), .I1(n4684), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8293.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8294 (.I0(\i14/fifo_inst/buff[116][2] ), .I1(\i14/fifo_inst/buff[118][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8294.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8295 (.I0(\i14/fifo_inst/buff[119][2] ), .I1(\i14/fifo_inst/buff[117][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8295.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8296 (.I0(n4687), .I1(n4688), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8296.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8297 (.I0(\i14/fifo_inst/buff[124][2] ), .I1(\i14/fifo_inst/buff[126][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8297.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8298 (.I0(\i14/fifo_inst/buff[127][2] ), .I1(\i14/fifo_inst/buff[125][2] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8298.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8299 (.I0(n4690), .I1(n4691), .I2(n4364), .O(n4692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8299.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8300 (.I0(\i14/fifo_inst/buff[120][2] ), .I1(\i14/fifo_inst/buff[122][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8300.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8301 (.I0(\i14/fifo_inst/buff[123][2] ), .I1(\i14/fifo_inst/buff[121][2] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8301.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8302 (.I0(n4694), .I1(n4693), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8302.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8303 (.I0(n4686), .I1(n4689), .I2(n4692), .I3(n4695), 
            .O(n4696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8303.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8304 (.I0(n4696), .I1(n4683), .I2(n4372), .I3(n4373), 
            .O(n4697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8304.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8305 (.I0(n4588), .I1(n4670), .I2(n4697), .I3(n4416), 
            .O(n4698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8305.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8306 (.I0(n4471), .I1(n4588), .I2(n4643), .I3(n4698), 
            .O(\fifo_inst/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__8306.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__8307 (.I0(\i14/fifo_inst/buff[20][3] ), .I1(\i14/fifo_inst/buff[22][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4699)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8307.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8308 (.I0(\i14/fifo_inst/buff[23][3] ), .I1(\i14/fifo_inst/buff[21][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4700)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8308.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8309 (.I0(n4699), .I1(n4700), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8309.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8310 (.I0(\i14/fifo_inst/buff[16][3] ), .I1(\i14/fifo_inst/buff[18][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4702)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8310.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8311 (.I0(\i14/fifo_inst/buff[19][3] ), .I1(\i14/fifo_inst/buff[17][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8311.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8312 (.I0(n4703), .I1(n4702), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8312.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8313 (.I0(\i14/fifo_inst/buff[24][3] ), .I1(\i14/fifo_inst/buff[26][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8313.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8314 (.I0(\i14/fifo_inst/buff[27][3] ), .I1(\i14/fifo_inst/buff[25][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8314.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8315 (.I0(n4358), .I1(n4705), .I2(n4706), .O(n4707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8315.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8316 (.I0(\i14/fifo_inst/buff[28][3] ), .I1(\i14/fifo_inst/buff[30][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8316.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8317 (.I0(\i14/fifo_inst/buff[31][3] ), .I1(\i14/fifo_inst/buff[29][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8317.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8318 (.I0(n4709), .I1(n4708), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4364), .O(n4710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8318.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8319 (.I0(n4701), .I1(n4704), .I2(n4707), .I3(n4710), 
            .O(n4711)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8319.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8320 (.I0(\i14/fifo_inst/buff[4][3] ), .I1(\i14/fifo_inst/buff[6][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4712)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8320.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8321 (.I0(\i14/fifo_inst/buff[7][3] ), .I1(\i14/fifo_inst/buff[5][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8321.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8322 (.I0(n4712), .I1(n4713), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8322.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8323 (.I0(\i14/fifo_inst/buff[8][3] ), .I1(\i14/fifo_inst/buff[10][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8323.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8324 (.I0(\i14/fifo_inst/buff[11][3] ), .I1(\i14/fifo_inst/buff[9][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8324.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8325 (.I0(n4716), .I1(n4715), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8325.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8326 (.I0(\i14/fifo_inst/buff[12][3] ), .I1(\i14/fifo_inst/buff[14][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8326.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8327 (.I0(\i14/fifo_inst/buff[15][3] ), .I1(\i14/fifo_inst/buff[13][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8327.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8328 (.I0(n4718), .I1(n4719), .I2(n4364), .O(n4720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8328.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8329 (.I0(\i14/fifo_inst/buff[0][3] ), .I1(\i14/fifo_inst/buff[2][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8329.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8330 (.I0(\i14/fifo_inst/buff[3][3] ), .I1(\i14/fifo_inst/buff[1][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8330.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8331 (.I0(n4368), .I1(n4721), .I2(n4722), .O(n4723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8331.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8332 (.I0(n4714), .I1(n4717), .I2(n4720), .I3(n4723), 
            .O(n4724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8332.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8333 (.I0(n4724), .I1(n4711), .I2(n4372), .I3(n4373), 
            .O(n4725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8333.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8334 (.I0(\i14/fifo_inst/buff[52][3] ), .I1(\i14/fifo_inst/buff[54][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4726)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8334.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8335 (.I0(\i14/fifo_inst/buff[55][3] ), .I1(\i14/fifo_inst/buff[53][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8335.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8336 (.I0(n4726), .I1(n4727), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8336.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8337 (.I0(\i14/fifo_inst/buff[56][3] ), .I1(\i14/fifo_inst/buff[58][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8337.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8338 (.I0(\i14/fifo_inst/buff[59][3] ), .I1(\i14/fifo_inst/buff[57][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4730)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8338.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8339 (.I0(n4730), .I1(n4729), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8339.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8340 (.I0(\i14/fifo_inst/buff[60][3] ), .I1(\i14/fifo_inst/buff[62][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8340.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8341 (.I0(\i14/fifo_inst/buff[63][3] ), .I1(\i14/fifo_inst/buff[61][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8341.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8342 (.I0(n4732), .I1(n4733), .I2(n4364), .O(n4734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8342.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8343 (.I0(\i14/fifo_inst/buff[48][3] ), .I1(\i14/fifo_inst/buff[50][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8343.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8344 (.I0(\i14/fifo_inst/buff[51][3] ), .I1(\i14/fifo_inst/buff[49][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8344.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8345 (.I0(n4368), .I1(n4735), .I2(n4736), .O(n4737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8345.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8346 (.I0(n4728), .I1(n4731), .I2(n4734), .I3(n4737), 
            .O(n4738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8346.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8347 (.I0(\i14/fifo_inst/buff[32][3] ), .I1(\i14/fifo_inst/buff[34][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8347.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8348 (.I0(\i14/fifo_inst/buff[35][3] ), .I1(\i14/fifo_inst/buff[33][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8348.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8349 (.I0(n4368), .I1(n4739), .I2(n4740), .O(n4741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8349.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8350 (.I0(\i14/fifo_inst/buff[40][3] ), .I1(\i14/fifo_inst/buff[42][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8350.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8351 (.I0(\i14/fifo_inst/buff[43][3] ), .I1(\i14/fifo_inst/buff[41][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8351.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8352 (.I0(n4743), .I1(n4742), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8352.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8353 (.I0(\i14/fifo_inst/buff[44][3] ), .I1(\i14/fifo_inst/buff[46][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8353.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8354 (.I0(\i14/fifo_inst/buff[47][3] ), .I1(\i14/fifo_inst/buff[45][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8354.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8355 (.I0(n4746), .I1(n4745), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4364), .O(n4747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8355.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8356 (.I0(\i14/fifo_inst/buff[36][3] ), .I1(\i14/fifo_inst/buff[38][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8356.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8357 (.I0(\i14/fifo_inst/buff[39][3] ), .I1(\i14/fifo_inst/buff[37][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8357.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8358 (.I0(n4748), .I1(n4749), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8358.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8359 (.I0(n4741), .I1(n4744), .I2(n4747), .I3(n4750), 
            .O(n4751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8359.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8360 (.I0(n4751), .I1(n4738), .I2(n4372), .I3(n4725), 
            .O(n4752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3f50 */ ;
    defparam LUT__8360.LUTMASK = 16'h3f50;
    EFX_LUT4 LUT__8361 (.I0(\i14/fifo_inst/buff[112][3] ), .I1(\i14/fifo_inst/buff[114][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8361.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8362 (.I0(\i14/fifo_inst/buff[115][3] ), .I1(\i14/fifo_inst/buff[113][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8362.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8363 (.I0(n4754), .I1(n4753), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8363.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8364 (.I0(\i14/fifo_inst/buff[124][3] ), .I1(\i14/fifo_inst/buff[126][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8364.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8365 (.I0(\i14/fifo_inst/buff[127][3] ), .I1(\i14/fifo_inst/buff[125][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8365.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8366 (.I0(n4757), .I1(n4756), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4364), .O(n4758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8366.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8367 (.I0(\i14/fifo_inst/buff[116][3] ), .I1(\i14/fifo_inst/buff[118][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8367.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8368 (.I0(\i14/fifo_inst/buff[119][3] ), .I1(\i14/fifo_inst/buff[117][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8368.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8369 (.I0(n4759), .I1(n4760), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8369.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8370 (.I0(\i14/fifo_inst/buff[120][3] ), .I1(\i14/fifo_inst/buff[122][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8370.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8371 (.I0(\i14/fifo_inst/buff[123][3] ), .I1(\i14/fifo_inst/buff[121][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8371.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8372 (.I0(n4763), .I1(n4762), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8372.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8373 (.I0(n4755), .I1(n4758), .I2(n4761), .I3(n4764), 
            .O(n4765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8373.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8374 (.I0(\i14/fifo_inst/buff[91][3] ), .I1(\i14/fifo_inst/buff[89][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4766)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8374.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8375 (.I0(\i14/fifo_inst/buff[88][3] ), .I1(\i14/fifo_inst/buff[90][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8375.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8376 (.I0(n4767), .I1(n4766), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8376.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8377 (.I0(\i14/fifo_inst/buff[87][3] ), .I1(\i14/fifo_inst/buff[85][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8377.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8378 (.I0(\i14/fifo_inst/buff[84][3] ), .I1(\i14/fifo_inst/buff[86][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8378.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8379 (.I0(n4769), .I1(n4770), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8379.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8380 (.I0(\i14/fifo_inst/buff[80][3] ), .I1(\i14/fifo_inst/buff[82][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8380.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8381 (.I0(\i14/fifo_inst/buff[83][3] ), .I1(\i14/fifo_inst/buff[81][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8381.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8382 (.I0(n4773), .I1(n4772), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8382.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8383 (.I0(\i14/fifo_inst/buff[92][3] ), .I1(\i14/fifo_inst/buff[94][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8383.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8384 (.I0(\i14/fifo_inst/buff[95][3] ), .I1(\i14/fifo_inst/buff[93][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8384.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8385 (.I0(n4776), .I1(n4775), .I2(n4364), .I3(\fifo_inst/rd_index[5] ), 
            .O(n4777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8385.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8386 (.I0(n4768), .I1(n4771), .I2(n4774), .I3(n4777), 
            .O(n4778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8386.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8387 (.I0(n4765), .I1(n4372), .I2(n4778), .I3(n4373), 
            .O(n4779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__8387.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__8388 (.I0(\i14/fifo_inst/buff[72][3] ), .I1(\i14/fifo_inst/buff[74][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8388.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8389 (.I0(\i14/fifo_inst/buff[75][3] ), .I1(\i14/fifo_inst/buff[73][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8389.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8390 (.I0(n4781), .I1(n4780), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8390.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8391 (.I0(\i14/fifo_inst/buff[68][3] ), .I1(\i14/fifo_inst/buff[70][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8391.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8392 (.I0(\i14/fifo_inst/buff[71][3] ), .I1(\i14/fifo_inst/buff[69][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8392.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8393 (.I0(n4783), .I1(n4784), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8393.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8394 (.I0(\i14/fifo_inst/buff[76][3] ), .I1(\i14/fifo_inst/buff[78][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8394.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8395 (.I0(\i14/fifo_inst/buff[79][3] ), .I1(\i14/fifo_inst/buff[77][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8395.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8396 (.I0(n4786), .I1(n4787), .I2(n4364), .O(n4788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8396.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8397 (.I0(\i14/fifo_inst/buff[64][3] ), .I1(\i14/fifo_inst/buff[66][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8397.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8398 (.I0(\i14/fifo_inst/buff[67][3] ), .I1(\i14/fifo_inst/buff[65][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8398.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8399 (.I0(n4790), .I1(n4789), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8399.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8400 (.I0(n4782), .I1(n4785), .I2(n4788), .I3(n4791), 
            .O(n4792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8400.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8401 (.I0(\i14/fifo_inst/buff[108][3] ), .I1(\i14/fifo_inst/buff[110][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8401.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8402 (.I0(\i14/fifo_inst/buff[111][3] ), .I1(\i14/fifo_inst/buff[109][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8402.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8403 (.I0(n4793), .I1(n4794), .I2(n4364), .O(n4795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8403.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8404 (.I0(\i14/fifo_inst/buff[96][3] ), .I1(\i14/fifo_inst/buff[98][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8404.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8405 (.I0(\i14/fifo_inst/buff[99][3] ), .I1(\i14/fifo_inst/buff[97][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8405.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8406 (.I0(n4368), .I1(n4796), .I2(n4797), .O(n4798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8406.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8407 (.I0(\i14/fifo_inst/buff[100][3] ), .I1(\i14/fifo_inst/buff[102][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8407.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8408 (.I0(\i14/fifo_inst/buff[103][3] ), .I1(\i14/fifo_inst/buff[101][3] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8408.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8409 (.I0(n4799), .I1(n4800), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8409.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8410 (.I0(\i14/fifo_inst/buff[104][3] ), .I1(\i14/fifo_inst/buff[106][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8410.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8411 (.I0(\i14/fifo_inst/buff[107][3] ), .I1(\i14/fifo_inst/buff[105][3] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8411.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8412 (.I0(n4803), .I1(n4802), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8412.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8413 (.I0(n4795), .I1(n4798), .I2(n4801), .I3(n4804), 
            .O(n4805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8413.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8414 (.I0(n4805), .I1(n4792), .I2(n4373), .I3(n4372), 
            .O(n4806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8414.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8415 (.I0(n4779), .I1(n4806), .I2(n4416), .I3(n4471), 
            .O(n4807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8415.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8416 (.I0(rx_en_fifo), .I1(n4319), .I2(\rx_d[3] ), .O(n4808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__8416.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__8417 (.I0(n4807), .I1(n4808), .I2(n4752), .I3(n4473), 
            .O(\fifo_inst/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__8417.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__8418 (.I0(rx_en_fifo), .I1(n4319), .O(n4809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8418.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8419 (.I0(\i14/fifo_inst/buff[8][4] ), .I1(\i14/fifo_inst/buff[10][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8419.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8420 (.I0(\i14/fifo_inst/buff[11][4] ), .I1(\i14/fifo_inst/buff[9][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8420.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8421 (.I0(n4811), .I1(n4810), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8421.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8422 (.I0(\i14/fifo_inst/buff[4][4] ), .I1(\i14/fifo_inst/buff[6][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8422.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8423 (.I0(\i14/fifo_inst/buff[7][4] ), .I1(\i14/fifo_inst/buff[5][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4814)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8423.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8424 (.I0(n4813), .I1(n4814), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n4815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8424.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8425 (.I0(\i14/fifo_inst/buff[12][4] ), .I1(\i14/fifo_inst/buff[14][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8425.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8426 (.I0(\i14/fifo_inst/buff[15][4] ), .I1(\i14/fifo_inst/buff[13][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8426.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8427 (.I0(\i14/fifo_inst/buff[3][4] ), .I1(\i14/fifo_inst/buff[1][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8427.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8428 (.I0(\i14/fifo_inst/buff[0][4] ), .I1(\i14/fifo_inst/buff[2][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8428.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8429 (.I0(n4819), .I1(n4818), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8429.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8430 (.I0(n4817), .I1(n4816), .I2(n4364), .I3(n4820), 
            .O(n4821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8430.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8431 (.I0(n4815), .I1(n4812), .I2(n4821), .I3(n4373), 
            .O(n4822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8431.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8432 (.I0(\i14/fifo_inst/buff[19][4] ), .I1(\i14/fifo_inst/buff[17][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8432.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8433 (.I0(\i14/fifo_inst/buff[16][4] ), .I1(\i14/fifo_inst/buff[18][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8433.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8434 (.I0(\i14/fifo_inst/buff[20][4] ), .I1(\i14/fifo_inst/buff[22][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8434.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8435 (.I0(\i14/fifo_inst/buff[23][4] ), .I1(\i14/fifo_inst/buff[21][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8435.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8436 (.I0(n4825), .I1(n4826), .I2(n4355), .I3(n4475), 
            .O(n4827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8436.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8437 (.I0(n4824), .I1(n4355), .I2(n4823), .I3(n4827), 
            .O(n4828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8437.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8438 (.I0(\i14/fifo_inst/buff[27][4] ), .I1(\i14/fifo_inst/buff[25][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8438.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8439 (.I0(\i14/fifo_inst/buff[24][4] ), .I1(\i14/fifo_inst/buff[26][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8439.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8440 (.I0(\i14/fifo_inst/buff[31][4] ), .I1(\i14/fifo_inst/buff[29][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8440.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8441 (.I0(\i14/fifo_inst/buff[28][4] ), .I1(\i14/fifo_inst/buff[30][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8441.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8442 (.I0(n4831), .I1(n4832), .I2(n4355), .I3(n4475), 
            .O(n4833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8442.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8443 (.I0(n4830), .I1(n4355), .I2(n4829), .I3(n4833), 
            .O(n4834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8443.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8444 (.I0(n4371), .I1(\fifo_inst/rd_index[4] ), .I2(\fifo_inst/rd_index[5] ), 
            .I3(\fifo_inst/rd_index[6] ), .O(n4835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ff8 */ ;
    defparam LUT__8444.LUTMASK = 16'h7ff8;
    EFX_LUT4 LUT__8445 (.I0(n4834), .I1(n4828), .I2(n4373), .I3(n4835), 
            .O(n4836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8445.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8446 (.I0(\i14/fifo_inst/buff[80][4] ), .I1(\i14/fifo_inst/buff[81][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haffc */ ;
    defparam LUT__8446.LUTMASK = 16'haffc;
    EFX_LUT4 LUT__8447 (.I0(\i14/fifo_inst/buff[82][4] ), .I1(\i14/fifo_inst/buff[83][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfacf */ ;
    defparam LUT__8447.LUTMASK = 16'hfacf;
    EFX_LUT4 LUT__8448 (.I0(\i14/fifo_inst/buff[88][4] ), .I1(\i14/fifo_inst/buff[90][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8448.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8449 (.I0(\i14/fifo_inst/buff[91][4] ), .I1(\i14/fifo_inst/buff[89][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n4839), .O(n4840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8449.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8450 (.I0(n4838), .I1(n4837), .I2(n4840), .I3(n4475), 
            .O(n4841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__8450.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__8451 (.I0(\i14/fifo_inst/buff[84][4] ), .I1(\i14/fifo_inst/buff[86][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8451.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8452 (.I0(\i14/fifo_inst/buff[87][4] ), .I1(\i14/fifo_inst/buff[85][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8452.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8453 (.I0(\i14/fifo_inst/buff[92][4] ), .I1(\i14/fifo_inst/buff[94][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8453.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8454 (.I0(\i14/fifo_inst/buff[95][4] ), .I1(\i14/fifo_inst/buff[93][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n4844), .O(n4845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8454.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8455 (.I0(n4843), .I1(n4842), .I2(n4845), .I3(n4475), 
            .O(n4846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__8455.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__8456 (.I0(rx_en_fifo_length), .I1(n4352), .I2(n4319), 
            .I3(n4373), .O(n4847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8456.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8457 (.I0(n4846), .I1(n4841), .I2(n4355), .I3(n4847), 
            .O(n4848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8457.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8458 (.I0(\i14/fifo_inst/buff[64][4] ), .I1(\i14/fifo_inst/buff[66][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8458.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8459 (.I0(\i14/fifo_inst/buff[65][4] ), .I1(\i14/fifo_inst/buff[67][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n4849), .O(n4850)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__8459.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__8460 (.I0(\i14/fifo_inst/buff[68][4] ), .I1(\i14/fifo_inst/buff[70][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8460.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8461 (.I0(\i14/fifo_inst/buff[71][4] ), .I1(\i14/fifo_inst/buff[69][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n4851), .O(n4852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8461.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8462 (.I0(n4852), .I1(n4850), .I2(n4355), .I3(n4475), 
            .O(n4853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha300 */ ;
    defparam LUT__8462.LUTMASK = 16'ha300;
    EFX_LUT4 LUT__8463 (.I0(n4371), .I1(\fifo_inst/rd_index[4] ), .I2(\fifo_inst/rd_index[6] ), 
            .I3(\fifo_inst/rd_index[5] ), .O(n4854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf78f */ ;
    defparam LUT__8463.LUTMASK = 16'hf78f;
    EFX_LUT4 LUT__8464 (.I0(rx_en_fifo_length), .I1(n4352), .I2(n4319), 
            .I3(n4854), .O(n4855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8464.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8465 (.I0(\i14/fifo_inst/buff[72][4] ), .I1(\i14/fifo_inst/buff[73][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haffc */ ;
    defparam LUT__8465.LUTMASK = 16'haffc;
    EFX_LUT4 LUT__8466 (.I0(\i14/fifo_inst/buff[74][4] ), .I1(\i14/fifo_inst/buff[75][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfacf */ ;
    defparam LUT__8466.LUTMASK = 16'hfacf;
    EFX_LUT4 LUT__8467 (.I0(\i14/fifo_inst/buff[76][4] ), .I1(\i14/fifo_inst/buff[78][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8467.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8468 (.I0(\i14/fifo_inst/buff[79][4] ), .I1(\i14/fifo_inst/buff[77][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8468.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8469 (.I0(n4858), .I1(n4859), .I2(n4355), .I3(n4475), 
            .O(n4860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8469.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8470 (.I0(n4355), .I1(n4857), .I2(n4856), .I3(n4860), 
            .O(n4861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__8470.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__8471 (.I0(rx_en_fifo_length), .I1(n4352), .I2(n4319), 
            .I3(n4373), .O(n4862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8471.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8472 (.I0(n4853), .I1(n4861), .I2(n4862), .I3(n4855), 
            .O(n4863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8472.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8473 (.I0(n4848), .I1(n4863), .I2(n4822), .I3(n4836), 
            .O(n4864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__8473.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__8474 (.I0(\i14/fifo_inst/buff[108][4] ), .I1(\i14/fifo_inst/buff[110][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8474.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8475 (.I0(\i14/fifo_inst/buff[111][4] ), .I1(\i14/fifo_inst/buff[109][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8475.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8476 (.I0(\i14/fifo_inst/buff[104][4] ), .I1(\i14/fifo_inst/buff[106][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8476.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8477 (.I0(\i14/fifo_inst/buff[107][4] ), .I1(\i14/fifo_inst/buff[105][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n4867), .O(n4868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8477.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8478 (.I0(n4866), .I1(n4865), .I2(n4868), .I3(n4355), 
            .O(n4869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__8478.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__8479 (.I0(\i14/fifo_inst/buff[99][4] ), .I1(\i14/fifo_inst/buff[97][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8479.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8480 (.I0(\i14/fifo_inst/buff[96][4] ), .I1(\i14/fifo_inst/buff[98][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8480.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8481 (.I0(\i14/fifo_inst/buff[100][4] ), .I1(\i14/fifo_inst/buff[102][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8481.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8482 (.I0(\i14/fifo_inst/buff[103][4] ), .I1(\i14/fifo_inst/buff[101][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n4872), .O(n4873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8482.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8483 (.I0(n4871), .I1(n4870), .I2(n4873), .I3(n4355), 
            .O(n4874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__8483.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__8484 (.I0(n4874), .I1(n4869), .I2(n4373), .I3(n4475), 
            .O(n4875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8484.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8485 (.I0(\i14/fifo_inst/buff[116][4] ), .I1(\i14/fifo_inst/buff[118][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8485.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8486 (.I0(\i14/fifo_inst/buff[119][4] ), .I1(\i14/fifo_inst/buff[117][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8486.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8487 (.I0(\i14/fifo_inst/buff[112][4] ), .I1(\i14/fifo_inst/buff[114][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8487.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8488 (.I0(\i14/fifo_inst/buff[115][4] ), .I1(\i14/fifo_inst/buff[113][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8488.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8489 (.I0(n4879), .I1(n4355), .I2(n4878), .I3(n4475), 
            .O(n4880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8489.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8490 (.I0(n4876), .I1(n4877), .I2(n4355), .I3(n4880), 
            .O(n4881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8490.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8491 (.I0(\i14/fifo_inst/buff[124][4] ), .I1(\i14/fifo_inst/buff[126][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8491.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8492 (.I0(\i14/fifo_inst/buff[127][4] ), .I1(\i14/fifo_inst/buff[125][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8492.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8493 (.I0(\i14/fifo_inst/buff[120][4] ), .I1(\i14/fifo_inst/buff[122][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8493.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8494 (.I0(\i14/fifo_inst/buff[123][4] ), .I1(\i14/fifo_inst/buff[121][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8494.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8495 (.I0(n4885), .I1(n4355), .I2(n4884), .I3(n4475), 
            .O(n4886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8495.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8496 (.I0(n4882), .I1(n4883), .I2(n4355), .I3(n4886), 
            .O(n4887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8496.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8497 (.I0(n4372), .I1(\fifo_inst/rd_index[6] ), .O(n4888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8497.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8498 (.I0(n4887), .I1(n4881), .I2(n4373), .I3(n4888), 
            .O(n4889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8498.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8499 (.I0(\i14/fifo_inst/buff[43][4] ), .I1(\i14/fifo_inst/buff[41][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8499.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8500 (.I0(\i14/fifo_inst/buff[40][4] ), .I1(\i14/fifo_inst/buff[42][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8500.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8501 (.I0(\i14/fifo_inst/buff[44][4] ), .I1(\i14/fifo_inst/buff[46][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8501.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8502 (.I0(\i14/fifo_inst/buff[47][4] ), .I1(\i14/fifo_inst/buff[45][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n4892), .O(n4893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8502.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8503 (.I0(n4891), .I1(n4890), .I2(n4893), .I3(n4355), 
            .O(n4894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__8503.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__8504 (.I0(\i14/fifo_inst/buff[35][4] ), .I1(\i14/fifo_inst/buff[33][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8504.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8505 (.I0(\i14/fifo_inst/buff[32][4] ), .I1(\i14/fifo_inst/buff[34][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8505.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8506 (.I0(\i14/fifo_inst/buff[36][4] ), .I1(\i14/fifo_inst/buff[38][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8506.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8507 (.I0(\i14/fifo_inst/buff[39][4] ), .I1(\i14/fifo_inst/buff[37][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n4897), .O(n4898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8507.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8508 (.I0(n4896), .I1(n4895), .I2(n4898), .I3(n4355), 
            .O(n4899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__8508.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__8509 (.I0(n4899), .I1(n4894), .I2(n4373), .I3(n4475), 
            .O(n4900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8509.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8510 (.I0(\i14/fifo_inst/buff[60][4] ), .I1(\i14/fifo_inst/buff[62][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8510.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8511 (.I0(\i14/fifo_inst/buff[63][4] ), .I1(\i14/fifo_inst/buff[61][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8511.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8512 (.I0(\i14/fifo_inst/buff[59][4] ), .I1(\i14/fifo_inst/buff[57][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8512.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8513 (.I0(\i14/fifo_inst/buff[56][4] ), .I1(\i14/fifo_inst/buff[58][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8513.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8514 (.I0(n4904), .I1(n4355), .I2(n4903), .I3(n4475), 
            .O(n4905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8514.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8515 (.I0(n4901), .I1(n4902), .I2(n4355), .I3(n4905), 
            .O(n4906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8515.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8516 (.I0(\i14/fifo_inst/buff[52][4] ), .I1(\i14/fifo_inst/buff[54][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8516.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8517 (.I0(\i14/fifo_inst/buff[55][4] ), .I1(\i14/fifo_inst/buff[53][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8517.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8518 (.I0(\i14/fifo_inst/buff[51][4] ), .I1(\i14/fifo_inst/buff[49][4] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8518.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8519 (.I0(\i14/fifo_inst/buff[48][4] ), .I1(\i14/fifo_inst/buff[50][4] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8519.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8520 (.I0(n4910), .I1(n4355), .I2(n4909), .I3(n4475), 
            .O(n4911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8520.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8521 (.I0(n4907), .I1(n4908), .I2(n4355), .I3(n4911), 
            .O(n4912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8521.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8522 (.I0(\fifo_inst/rd_index[6] ), .I1(n4372), .O(n4913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8522.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8523 (.I0(n4912), .I1(n4906), .I2(n4373), .I3(n4913), 
            .O(n4914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8523.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8524 (.I0(n4900), .I1(n4914), .I2(n4875), .I3(n4889), 
            .O(n4915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__8524.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__8525 (.I0(n4864), .I1(n4915), .I2(n4809), .I3(\rx_d[4] ), 
            .O(\fifo_inst/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888 */ ;
    defparam LUT__8525.LUTMASK = 16'hf888;
    EFX_LUT4 LUT__8526 (.I0(\i14/fifo_inst/buff[0][5] ), .I1(\i14/fifo_inst/buff[2][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8526.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8527 (.I0(\i14/fifo_inst/buff[3][5] ), .I1(\i14/fifo_inst/buff[1][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8527.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8528 (.I0(n4917), .I1(n4916), .I2(n4355), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8528.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8529 (.I0(\i14/fifo_inst/buff[7][5] ), .I1(\i14/fifo_inst/buff[5][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8529.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8530 (.I0(\i14/fifo_inst/buff[4][5] ), .I1(\i14/fifo_inst/buff[6][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8530.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8531 (.I0(n4920), .I1(n4919), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4355), .O(n4921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8531.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8532 (.I0(n4921), .I1(n4918), .I2(n4475), .I3(n4373), 
            .O(n4922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8532.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8533 (.I0(\i14/fifo_inst/buff[12][5] ), .I1(\i14/fifo_inst/buff[14][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8533.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8534 (.I0(\i14/fifo_inst/buff[15][5] ), .I1(\i14/fifo_inst/buff[13][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8534.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8535 (.I0(n4924), .I1(n4923), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4355), .O(n4925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8535.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8536 (.I0(\fifo_inst/rd_index[0] ), .I1(\fifo_inst/rd_index[1] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(\i14/fifo_inst/buff[8][5] ), 
            .O(n4926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8536.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8537 (.I0(\i14/fifo_inst/buff[9][5] ), .I1(\i14/fifo_inst/buff[11][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8537.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8538 (.I0(\i14/fifo_inst/buff[10][5] ), .I1(\fifo_inst/rd_index[0] ), 
            .I2(\fifo_inst/rd_index[2] ), .I3(n4927), .O(n4928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__8538.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__8539 (.I0(n4925), .I1(n4926), .I2(n4475), .I3(n4928), 
            .O(n4929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8539.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8540 (.I0(\i14/fifo_inst/buff[28][5] ), .I1(\i14/fifo_inst/buff[30][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8540.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8541 (.I0(\i14/fifo_inst/buff[31][5] ), .I1(\i14/fifo_inst/buff[29][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8541.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8542 (.I0(\i14/fifo_inst/buff[24][5] ), .I1(\i14/fifo_inst/buff[26][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8542.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8543 (.I0(\i14/fifo_inst/buff[27][5] ), .I1(\i14/fifo_inst/buff[25][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8543.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8544 (.I0(n4933), .I1(n4355), .I2(n4932), .I3(n4475), 
            .O(n4934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8544.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8545 (.I0(n4930), .I1(n4931), .I2(n4355), .I3(n4934), 
            .O(n4935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8545.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8546 (.I0(\i14/fifo_inst/buff[16][5] ), .I1(\i14/fifo_inst/buff[18][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8546.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8547 (.I0(\i14/fifo_inst/buff[19][5] ), .I1(\i14/fifo_inst/buff[17][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8547.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8548 (.I0(\i14/fifo_inst/buff[20][5] ), .I1(\i14/fifo_inst/buff[21][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haffc */ ;
    defparam LUT__8548.LUTMASK = 16'haffc;
    EFX_LUT4 LUT__8549 (.I0(\i14/fifo_inst/buff[22][5] ), .I1(\i14/fifo_inst/buff[23][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfacf */ ;
    defparam LUT__8549.LUTMASK = 16'hfacf;
    EFX_LUT4 LUT__8550 (.I0(n4938), .I1(n4939), .I2(n4355), .I3(n4475), 
            .O(n4940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__8550.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__8551 (.I0(n4937), .I1(n4355), .I2(n4936), .I3(n4940), 
            .O(n4941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8551.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8552 (.I0(n4935), .I1(n4941), .I2(n4373), .O(n4942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8552.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8553 (.I0(n4929), .I1(n4922), .I2(n4942), .I3(n4835), 
            .O(n4943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__8553.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__8554 (.I0(\i14/fifo_inst/buff[107][5] ), .I1(\i14/fifo_inst/buff[105][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8554.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8555 (.I0(\i14/fifo_inst/buff[104][5] ), .I1(\i14/fifo_inst/buff[106][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8555.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8556 (.I0(n4945), .I1(n4355), .I2(n4944), .I3(n4475), 
            .O(n4946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8556.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8557 (.I0(\i14/fifo_inst/buff[111][5] ), .I1(\i14/fifo_inst/buff[109][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8557.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8558 (.I0(\i14/fifo_inst/buff[108][5] ), .I1(\i14/fifo_inst/buff[110][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8558.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8559 (.I0(n4948), .I1(n4947), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4355), .O(n4949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8559.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8560 (.I0(\i14/fifo_inst/buff[103][5] ), .I1(\i14/fifo_inst/buff[101][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8560.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8561 (.I0(\i14/fifo_inst/buff[100][5] ), .I1(\i14/fifo_inst/buff[102][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8561.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8562 (.I0(\i14/fifo_inst/buff[99][5] ), .I1(\i14/fifo_inst/buff[97][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8562.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8563 (.I0(\i14/fifo_inst/buff[96][5] ), .I1(\i14/fifo_inst/buff[98][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8563.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8564 (.I0(n4953), .I1(n4355), .I2(n4952), .I3(n4475), 
            .O(n4954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8564.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8565 (.I0(n4950), .I1(n4951), .I2(n4355), .I3(n4954), 
            .O(n4955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8565.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8566 (.I0(n4949), .I1(n4946), .I2(n4955), .I3(n4373), 
            .O(n4956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__8566.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__8567 (.I0(\i14/fifo_inst/buff[120][5] ), .I1(\i14/fifo_inst/buff[122][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8567.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8568 (.I0(\i14/fifo_inst/buff[123][5] ), .I1(\i14/fifo_inst/buff[121][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n4957), .O(n4958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8568.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8569 (.I0(\i14/fifo_inst/buff[124][5] ), .I1(\i14/fifo_inst/buff[126][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8569.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8570 (.I0(\i14/fifo_inst/buff[127][5] ), .I1(\i14/fifo_inst/buff[125][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n4959), .O(n4960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8570.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8571 (.I0(n4960), .I1(n4958), .I2(n4475), .I3(n4355), 
            .O(n4961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__8571.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__8572 (.I0(\i14/fifo_inst/buff[116][5] ), .I1(\i14/fifo_inst/buff[118][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8572.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8573 (.I0(\i14/fifo_inst/buff[119][5] ), .I1(\i14/fifo_inst/buff[117][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8573.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8574 (.I0(\i14/fifo_inst/buff[115][5] ), .I1(\i14/fifo_inst/buff[113][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8574.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8575 (.I0(\i14/fifo_inst/buff[112][5] ), .I1(\i14/fifo_inst/buff[114][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8575.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8576 (.I0(n4965), .I1(n4355), .I2(n4964), .I3(n4475), 
            .O(n4966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8576.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8577 (.I0(n4962), .I1(n4963), .I2(n4355), .I3(n4966), 
            .O(n4967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8577.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8578 (.I0(n4967), .I1(n4961), .I2(n4373), .I3(n4888), 
            .O(n4968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8578.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8579 (.I0(\i14/fifo_inst/buff[43][5] ), .I1(\i14/fifo_inst/buff[41][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8579.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8580 (.I0(\i14/fifo_inst/buff[40][5] ), .I1(\i14/fifo_inst/buff[42][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8580.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8581 (.I0(\i14/fifo_inst/buff[44][5] ), .I1(\i14/fifo_inst/buff[46][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8581.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8582 (.I0(\i14/fifo_inst/buff[47][5] ), .I1(\i14/fifo_inst/buff[45][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n4971), .O(n4972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8582.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8583 (.I0(n4970), .I1(n4969), .I2(n4972), .I3(n4355), 
            .O(n4973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__8583.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__8584 (.I0(\i14/fifo_inst/buff[35][5] ), .I1(\i14/fifo_inst/buff[33][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8584.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8585 (.I0(\i14/fifo_inst/buff[32][5] ), .I1(\i14/fifo_inst/buff[34][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8585.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8586 (.I0(\i14/fifo_inst/buff[36][5] ), .I1(\i14/fifo_inst/buff[38][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8586.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8587 (.I0(\i14/fifo_inst/buff[39][5] ), .I1(\i14/fifo_inst/buff[37][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n4976), .O(n4977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8587.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8588 (.I0(n4975), .I1(n4974), .I2(n4977), .I3(n4355), 
            .O(n4978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__8588.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__8589 (.I0(n4978), .I1(n4973), .I2(n4373), .I3(n4475), 
            .O(n4979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8589.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8590 (.I0(\i14/fifo_inst/buff[55][5] ), .I1(\i14/fifo_inst/buff[53][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8590.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8591 (.I0(\i14/fifo_inst/buff[52][5] ), .I1(\i14/fifo_inst/buff[54][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4981)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8591.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8592 (.I0(\i14/fifo_inst/buff[51][5] ), .I1(\i14/fifo_inst/buff[49][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8592.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8593 (.I0(\i14/fifo_inst/buff[48][5] ), .I1(\i14/fifo_inst/buff[50][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8593.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8594 (.I0(n4982), .I1(n4983), .I2(n4981), .I3(n4355), 
            .O(n4984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__8594.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__8595 (.I0(n4980), .I1(n4355), .I2(n4984), .I3(n4475), 
            .O(n4985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__8595.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__8596 (.I0(\i14/fifo_inst/buff[60][5] ), .I1(\i14/fifo_inst/buff[62][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8596.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8597 (.I0(\i14/fifo_inst/buff[63][5] ), .I1(\i14/fifo_inst/buff[61][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8597.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8598 (.I0(\i14/fifo_inst/buff[59][5] ), .I1(\i14/fifo_inst/buff[57][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8598.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8599 (.I0(\i14/fifo_inst/buff[56][5] ), .I1(\i14/fifo_inst/buff[58][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8599.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8600 (.I0(n4989), .I1(n4355), .I2(n4988), .I3(n4475), 
            .O(n4990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8600.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8601 (.I0(n4986), .I1(n4987), .I2(n4355), .I3(n4990), 
            .O(n4991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8601.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8602 (.I0(n4985), .I1(n4991), .I2(n4373), .I3(n4913), 
            .O(n4992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8602.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8603 (.I0(n4979), .I1(n4992), .I2(n4956), .I3(n4968), 
            .O(n4993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__8603.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__8604 (.I0(\i14/fifo_inst/buff[92][5] ), .I1(\i14/fifo_inst/buff[94][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8604.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8605 (.I0(\i14/fifo_inst/buff[95][5] ), .I1(\i14/fifo_inst/buff[93][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n4995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8605.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8606 (.I0(n4994), .I1(n4995), .I2(n4355), .I3(n4475), 
            .O(n4996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8606.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8607 (.I0(\i14/fifo_inst/buff[91][5] ), .I1(\i14/fifo_inst/buff[89][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8607.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8608 (.I0(\i14/fifo_inst/buff[88][5] ), .I1(\i14/fifo_inst/buff[90][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n4998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8608.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8609 (.I0(n4998), .I1(n4997), .I2(n4355), .I3(\fifo_inst/rd_index[0] ), 
            .O(n4999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8609.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8610 (.I0(\i14/fifo_inst/buff[84][5] ), .I1(\i14/fifo_inst/buff[86][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8610.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8611 (.I0(\i14/fifo_inst/buff[87][5] ), .I1(\i14/fifo_inst/buff[85][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8611.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8612 (.I0(\i14/fifo_inst/buff[80][5] ), .I1(\i14/fifo_inst/buff[83][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8612.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8613 (.I0(\i14/fifo_inst/buff[82][5] ), .I1(\i14/fifo_inst/buff[81][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8613.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8614 (.I0(n5003), .I1(n4355), .I2(n5002), .I3(n4475), 
            .O(n5004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8614.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8615 (.I0(n5000), .I1(n5001), .I2(n4355), .I3(n5004), 
            .O(n5005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8615.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8616 (.I0(n4999), .I1(n4996), .I2(n5005), .I3(n4373), 
            .O(n5006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__8616.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__8617 (.I0(\i14/fifo_inst/buff[72][5] ), .I1(\i14/fifo_inst/buff[74][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n5007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8617.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8618 (.I0(\i14/fifo_inst/buff[75][5] ), .I1(\i14/fifo_inst/buff[73][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n5008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8618.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8619 (.I0(n5008), .I1(n5007), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8619.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8620 (.I0(\i14/fifo_inst/buff[64][5] ), .I1(\i14/fifo_inst/buff[66][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n5010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8620.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8621 (.I0(\i14/fifo_inst/buff[67][5] ), .I1(\i14/fifo_inst/buff[65][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n5011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8621.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8622 (.I0(n5011), .I1(n5010), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8622.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8623 (.I0(\i14/fifo_inst/buff[76][5] ), .I1(\i14/fifo_inst/buff[78][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8623.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8624 (.I0(\i14/fifo_inst/buff[79][5] ), .I1(\i14/fifo_inst/buff[77][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8624.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8625 (.I0(\i14/fifo_inst/buff[68][5] ), .I1(\i14/fifo_inst/buff[70][5] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8625.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8626 (.I0(\i14/fifo_inst/buff[71][5] ), .I1(\i14/fifo_inst/buff[69][5] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8626.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8627 (.I0(n5015), .I1(n5016), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n5017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8627.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8628 (.I0(n5014), .I1(n5013), .I2(n4364), .I3(n5017), 
            .O(n5018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8628.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8629 (.I0(n5012), .I1(n5009), .I2(n5018), .I3(n4373), 
            .O(n5019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8629.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8630 (.I0(n5019), .I1(n4854), .I2(n5006), .I3(n4471), 
            .O(n5020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8630.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8631 (.I0(n4809), .I1(\rx_d[5] ), .O(n5021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8631.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8632 (.I0(n4943), .I1(n5020), .I2(n4993), .I3(n5021), 
            .O(\fifo_inst/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40 */ ;
    defparam LUT__8632.LUTMASK = 16'hff40;
    EFX_LUT4 LUT__8633 (.I0(\i14/fifo_inst/buff[83][6] ), .I1(\i14/fifo_inst/buff[81][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8633.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8634 (.I0(\i14/fifo_inst/buff[80][6] ), .I1(\i14/fifo_inst/buff[82][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8634.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8635 (.I0(\i14/fifo_inst/buff[87][6] ), .I1(\i14/fifo_inst/buff[85][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8635.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8636 (.I0(n5022), .I1(n5023), .I2(n5024), .I3(n4355), 
            .O(n5025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__8636.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__8637 (.I0(n5025), .I1(n4475), .I2(n4373), .O(n5026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__8637.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__8638 (.I0(\i14/fifo_inst/buff[91][6] ), .I1(\i14/fifo_inst/buff[89][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8638.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8639 (.I0(\i14/fifo_inst/buff[88][6] ), .I1(\i14/fifo_inst/buff[90][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8639.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8640 (.I0(\i14/fifo_inst/buff[92][6] ), .I1(\i14/fifo_inst/buff[94][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8640.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8641 (.I0(\i14/fifo_inst/buff[95][6] ), .I1(\i14/fifo_inst/buff[93][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8641.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8642 (.I0(\i14/fifo_inst/buff[84][6] ), .I1(\i14/fifo_inst/buff[86][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8642.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8643 (.I0(n5029), .I1(n5030), .I2(n5031), .I3(n4475), 
            .O(n5032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__8643.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__8644 (.I0(n5027), .I1(n5028), .I2(n5032), .I3(n4355), 
            .O(n5033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__8644.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__8645 (.I0(n4355), .I1(n4475), .I2(n5033), .I3(n5026), 
            .O(n5034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc700 */ ;
    defparam LUT__8645.LUTMASK = 16'hc700;
    EFX_LUT4 LUT__8646 (.I0(\i14/fifo_inst/buff[64][6] ), .I1(\i14/fifo_inst/buff[66][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n5035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8646.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8647 (.I0(\i14/fifo_inst/buff[67][6] ), .I1(\i14/fifo_inst/buff[65][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n5036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8647.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8648 (.I0(n5036), .I1(n5035), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8648.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8649 (.I0(\i14/fifo_inst/buff[72][6] ), .I1(\i14/fifo_inst/buff[74][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n5038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8649.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8650 (.I0(\i14/fifo_inst/buff[75][6] ), .I1(\i14/fifo_inst/buff[73][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n5039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8650.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8651 (.I0(n5039), .I1(n5038), .I2(n4358), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8651.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8652 (.I0(\i14/fifo_inst/buff[68][6] ), .I1(\i14/fifo_inst/buff[70][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8652.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8653 (.I0(\i14/fifo_inst/buff[71][6] ), .I1(\i14/fifo_inst/buff[69][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8653.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8654 (.I0(n5041), .I1(n5042), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n5043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8654.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8655 (.I0(\i14/fifo_inst/buff[76][6] ), .I1(\i14/fifo_inst/buff[78][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n5044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8655.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8656 (.I0(\i14/fifo_inst/buff[79][6] ), .I1(\i14/fifo_inst/buff[77][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n5045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8656.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8657 (.I0(n5045), .I1(n5044), .I2(\fifo_inst/rd_index[0] ), 
            .I3(n4364), .O(n5046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8657.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8658 (.I0(n5037), .I1(n5040), .I2(n5043), .I3(n5046), 
            .O(n5047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8658.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8659 (.I0(n5047), .I1(n4373), .I2(n4854), .O(n5048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__8659.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__8660 (.I0(\i14/fifo_inst/buff[3][6] ), .I1(\i14/fifo_inst/buff[1][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8660.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8661 (.I0(\i14/fifo_inst/buff[2][6] ), .I1(\i14/fifo_inst/buff[0][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8661.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8662 (.I0(\i14/fifo_inst/buff[6][6] ), .I1(\i14/fifo_inst/buff[5][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8662.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8663 (.I0(\i14/fifo_inst/buff[4][6] ), .I1(\i14/fifo_inst/buff[7][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8663.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8664 (.I0(n5051), .I1(n5052), .I2(n4355), .I3(n4475), 
            .O(n5053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8664.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8665 (.I0(n5050), .I1(n4355), .I2(n5049), .I3(n5053), 
            .O(n5054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8665.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8666 (.I0(\i14/fifo_inst/buff[12][6] ), .I1(\i14/fifo_inst/buff[14][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8666.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8667 (.I0(\i14/fifo_inst/buff[15][6] ), .I1(\i14/fifo_inst/buff[13][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8667.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8668 (.I0(\i14/fifo_inst/buff[11][6] ), .I1(\i14/fifo_inst/buff[9][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8668.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8669 (.I0(\i14/fifo_inst/buff[8][6] ), .I1(\i14/fifo_inst/buff[10][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8669.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8670 (.I0(n5057), .I1(n5058), .I2(n5056), .I3(n4355), 
            .O(n5059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__8670.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__8671 (.I0(n5055), .I1(n4355), .I2(n4475), .I3(n5059), 
            .O(n5060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0c */ ;
    defparam LUT__8671.LUTMASK = 16'h0b0c;
    EFX_LUT4 LUT__8672 (.I0(n5054), .I1(n5060), .I2(n4862), .O(n5061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8672.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8673 (.I0(\i14/fifo_inst/buff[22][6] ), .I1(\i14/fifo_inst/buff[21][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8673.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8674 (.I0(\i14/fifo_inst/buff[20][6] ), .I1(\i14/fifo_inst/buff[23][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8674.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8675 (.I0(\i14/fifo_inst/buff[16][6] ), .I1(\i14/fifo_inst/buff[18][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8675.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8676 (.I0(\i14/fifo_inst/buff[19][6] ), .I1(\i14/fifo_inst/buff[17][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8676.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8677 (.I0(n5065), .I1(n4355), .I2(n5064), .I3(n4475), 
            .O(n5066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8677.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8678 (.I0(n5062), .I1(n5063), .I2(n4355), .I3(n5066), 
            .O(n5067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8678.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8679 (.I0(\i14/fifo_inst/buff[28][6] ), .I1(\i14/fifo_inst/buff[30][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8679.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8680 (.I0(\i14/fifo_inst/buff[31][6] ), .I1(\i14/fifo_inst/buff[29][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8680.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8681 (.I0(\i14/fifo_inst/buff[27][6] ), .I1(\i14/fifo_inst/buff[25][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8681.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8682 (.I0(\i14/fifo_inst/buff[24][6] ), .I1(\i14/fifo_inst/buff[26][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8682.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8683 (.I0(n5071), .I1(n4355), .I2(n5070), .I3(n4475), 
            .O(n5072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8683.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8684 (.I0(n5068), .I1(n5069), .I2(n4355), .I3(n5072), 
            .O(n5073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8684.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8685 (.I0(rx_en_fifo_length), .I1(n4352), .I2(n4319), 
            .I3(n4835), .O(n5074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8685.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8686 (.I0(n5073), .I1(n5067), .I2(n4847), .I3(n5074), 
            .O(n5075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8686.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8687 (.I0(n5061), .I1(n5075), .I2(n5034), .I3(n5048), 
            .O(n5076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__8687.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__8688 (.I0(\i14/fifo_inst/buff[123][6] ), .I1(\i14/fifo_inst/buff[121][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8688.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8689 (.I0(\i14/fifo_inst/buff[120][6] ), .I1(\i14/fifo_inst/buff[122][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8689.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8690 (.I0(\i14/fifo_inst/buff[124][6] ), .I1(\i14/fifo_inst/buff[126][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8690.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8691 (.I0(\i14/fifo_inst/buff[127][6] ), .I1(\i14/fifo_inst/buff[125][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8691.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8692 (.I0(n5079), .I1(n5080), .I2(n4355), .I3(n4475), 
            .O(n5081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8692.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8693 (.I0(n5078), .I1(n4355), .I2(n5077), .I3(n5081), 
            .O(n5082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8693.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8694 (.I0(\i14/fifo_inst/buff[115][6] ), .I1(\i14/fifo_inst/buff[113][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8694.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8695 (.I0(\i14/fifo_inst/buff[112][6] ), .I1(\i14/fifo_inst/buff[114][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8695.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8696 (.I0(\i14/fifo_inst/buff[116][6] ), .I1(\i14/fifo_inst/buff[118][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8696.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8697 (.I0(\i14/fifo_inst/buff[119][6] ), .I1(\i14/fifo_inst/buff[117][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8697.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8698 (.I0(n5085), .I1(n5086), .I2(n4355), .I3(n4475), 
            .O(n5087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8698.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8699 (.I0(n5084), .I1(n4355), .I2(n5083), .I3(n5087), 
            .O(n5088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8699.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8700 (.I0(n5082), .I1(n5088), .I2(n4373), .O(n5089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8700.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8701 (.I0(\i14/fifo_inst/buff[108][6] ), .I1(\i14/fifo_inst/buff[110][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8701.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8702 (.I0(\i14/fifo_inst/buff[111][6] ), .I1(\i14/fifo_inst/buff[109][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8702.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8703 (.I0(\i14/fifo_inst/buff[104][6] ), .I1(\i14/fifo_inst/buff[106][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8703.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8704 (.I0(\i14/fifo_inst/buff[107][6] ), .I1(\i14/fifo_inst/buff[105][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8704.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8705 (.I0(n5093), .I1(n4355), .I2(n5092), .I3(n4475), 
            .O(n5094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8705.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8706 (.I0(n5090), .I1(n5091), .I2(n4355), .I3(n5094), 
            .O(n5095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8706.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8707 (.I0(\i14/fifo_inst/buff[100][6] ), .I1(\i14/fifo_inst/buff[102][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8707.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8708 (.I0(\i14/fifo_inst/buff[103][6] ), .I1(\i14/fifo_inst/buff[101][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8708.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8709 (.I0(\i14/fifo_inst/buff[99][6] ), .I1(\i14/fifo_inst/buff[97][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8709.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8710 (.I0(\i14/fifo_inst/buff[96][6] ), .I1(\i14/fifo_inst/buff[98][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8710.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8711 (.I0(n5099), .I1(n4355), .I2(n5098), .I3(n4475), 
            .O(n5100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8711.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8712 (.I0(n5096), .I1(n5097), .I2(n4355), .I3(n5100), 
            .O(n5101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8712.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8713 (.I0(n5101), .I1(n4373), .I2(n5095), .I3(n4888), 
            .O(n5102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8713.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8714 (.I0(\i14/fifo_inst/buff[52][6] ), .I1(\i14/fifo_inst/buff[54][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8714.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8715 (.I0(\i14/fifo_inst/buff[55][6] ), .I1(\i14/fifo_inst/buff[53][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8715.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8716 (.I0(\i14/fifo_inst/buff[48][6] ), .I1(\i14/fifo_inst/buff[50][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8716.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8717 (.I0(\i14/fifo_inst/buff[51][6] ), .I1(\i14/fifo_inst/buff[49][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8717.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8718 (.I0(n5106), .I1(n4355), .I2(n5105), .I3(n4475), 
            .O(n5107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8718.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8719 (.I0(n5103), .I1(n5104), .I2(n4355), .I3(n5107), 
            .O(n5108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8719.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8720 (.I0(\i14/fifo_inst/buff[59][6] ), .I1(\i14/fifo_inst/buff[57][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8720.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8721 (.I0(\i14/fifo_inst/buff[56][6] ), .I1(\i14/fifo_inst/buff[58][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8721.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8722 (.I0(\i14/fifo_inst/buff[60][6] ), .I1(\i14/fifo_inst/buff[62][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8722.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8723 (.I0(\i14/fifo_inst/buff[63][6] ), .I1(\i14/fifo_inst/buff[61][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8723.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8724 (.I0(n5111), .I1(n5112), .I2(n4355), .I3(n4475), 
            .O(n5113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8724.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8725 (.I0(n5110), .I1(n4355), .I2(n5109), .I3(n5113), 
            .O(n5114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8725.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8726 (.I0(n5108), .I1(n5114), .I2(n4373), .O(n5115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8726.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8727 (.I0(\i14/fifo_inst/buff[35][6] ), .I1(\i14/fifo_inst/buff[33][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8727.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8728 (.I0(\i14/fifo_inst/buff[32][6] ), .I1(\i14/fifo_inst/buff[34][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8728.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8729 (.I0(\i14/fifo_inst/buff[36][6] ), .I1(\i14/fifo_inst/buff[38][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8729.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8730 (.I0(\i14/fifo_inst/buff[39][6] ), .I1(\i14/fifo_inst/buff[37][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8730.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8731 (.I0(n5118), .I1(n5119), .I2(n4355), .I3(n4475), 
            .O(n5120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8731.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8732 (.I0(n5117), .I1(n4355), .I2(n5116), .I3(n5120), 
            .O(n5121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8732.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8733 (.I0(\i14/fifo_inst/buff[44][6] ), .I1(\i14/fifo_inst/buff[46][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8733.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8734 (.I0(\i14/fifo_inst/buff[47][6] ), .I1(\i14/fifo_inst/buff[45][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8734.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8735 (.I0(\i14/fifo_inst/buff[40][6] ), .I1(\i14/fifo_inst/buff[42][6] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8735.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8736 (.I0(\i14/fifo_inst/buff[43][6] ), .I1(\i14/fifo_inst/buff[41][6] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8736.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8737 (.I0(n5125), .I1(n4355), .I2(n5124), .I3(n4475), 
            .O(n5126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8737.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8738 (.I0(n5122), .I1(n5123), .I2(n4355), .I3(n5126), 
            .O(n5127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8738.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8739 (.I0(n5127), .I1(n4373), .I2(n5121), .I3(n4913), 
            .O(n5128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8739.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8740 (.I0(n5115), .I1(n5128), .I2(n5089), .I3(n5102), 
            .O(n5129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__8740.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__8741 (.I0(n5076), .I1(n5129), .I2(n4809), .I3(\rx_d[6] ), 
            .O(\fifo_inst/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888 */ ;
    defparam LUT__8741.LUTMASK = 16'hf888;
    EFX_LUT4 LUT__8742 (.I0(\i14/fifo_inst/buff[3][7] ), .I1(\i14/fifo_inst/buff[1][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8742.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8743 (.I0(\i14/fifo_inst/buff[2][7] ), .I1(\i14/fifo_inst/buff[0][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8743.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8744 (.I0(\i14/fifo_inst/buff[7][7] ), .I1(\i14/fifo_inst/buff[5][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8744.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8745 (.I0(n5130), .I1(n5131), .I2(n5132), .I3(n4355), 
            .O(n5133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__8745.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__8746 (.I0(\i14/fifo_inst/buff[4][7] ), .I1(\i14/fifo_inst/buff[6][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8746.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8747 (.I0(\i14/fifo_inst/buff[12][7] ), .I1(\i14/fifo_inst/buff[14][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8747.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8748 (.I0(\i14/fifo_inst/buff[15][7] ), .I1(\i14/fifo_inst/buff[13][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8748.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8749 (.I0(n5135), .I1(n5136), .I2(n5134), .I3(n4475), 
            .O(n5137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__8749.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__8750 (.I0(\i14/fifo_inst/buff[11][7] ), .I1(\i14/fifo_inst/buff[9][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8750.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8751 (.I0(\i14/fifo_inst/buff[8][7] ), .I1(\i14/fifo_inst/buff[10][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8751.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8752 (.I0(n5138), .I1(n5139), .I2(n5137), .I3(n4355), 
            .O(n5140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__8752.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__8753 (.I0(n4355), .I1(n5133), .I2(n4475), .I3(n5140), 
            .O(n5141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h301f */ ;
    defparam LUT__8753.LUTMASK = 16'h301f;
    EFX_LUT4 LUT__8754 (.I0(\i14/fifo_inst/buff[20][7] ), .I1(\i14/fifo_inst/buff[22][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8754.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8755 (.I0(\i14/fifo_inst/buff[24][7] ), .I1(\i14/fifo_inst/buff[26][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8755.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8756 (.I0(\i14/fifo_inst/buff[27][7] ), .I1(\i14/fifo_inst/buff[25][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8756.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8757 (.I0(n5143), .I1(n5144), .I2(n5142), .I3(n4355), 
            .O(n5145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__8757.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__8758 (.I0(\i14/fifo_inst/buff[16][7] ), .I1(\i14/fifo_inst/buff[18][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8758.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8759 (.I0(\i14/fifo_inst/buff[19][7] ), .I1(\i14/fifo_inst/buff[17][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n5146), .O(n5147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8759.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8760 (.I0(n5147), .I1(n5145), .I2(n4355), .I3(n4475), 
            .O(n5148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h35f3 */ ;
    defparam LUT__8760.LUTMASK = 16'h35f3;
    EFX_LUT4 LUT__8761 (.I0(\i14/fifo_inst/buff[23][7] ), .I1(\i14/fifo_inst/buff[21][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8761.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8762 (.I0(\i14/fifo_inst/buff[28][7] ), .I1(\i14/fifo_inst/buff[30][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8762.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8763 (.I0(\i14/fifo_inst/buff[31][7] ), .I1(\i14/fifo_inst/buff[29][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8763.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8764 (.I0(n5150), .I1(n5151), .I2(n5149), .I3(n4475), 
            .O(n5152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__8764.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__8765 (.I0(n5152), .I1(n4355), .I2(n4847), .I3(n5148), 
            .O(n5153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__8765.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__8766 (.I0(n4862), .I1(n5141), .I2(n5074), .I3(n5153), 
            .O(n5154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__8766.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__8767 (.I0(\i14/fifo_inst/buff[72][7] ), .I1(\i14/fifo_inst/buff[74][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8767.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8768 (.I0(\i14/fifo_inst/buff[75][7] ), .I1(\i14/fifo_inst/buff[73][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n5155), .O(n5156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8768.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8769 (.I0(\i14/fifo_inst/buff[76][7] ), .I1(\i14/fifo_inst/buff[78][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8769.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8770 (.I0(\i14/fifo_inst/buff[79][7] ), .I1(\i14/fifo_inst/buff[77][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8770.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8771 (.I0(\i14/fifo_inst/buff[64][7] ), .I1(\i14/fifo_inst/buff[66][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n5159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8771.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8772 (.I0(\i14/fifo_inst/buff[67][7] ), .I1(\i14/fifo_inst/buff[65][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .O(n5160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8772.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8773 (.I0(n5160), .I1(n5159), .I2(n4368), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8773.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8774 (.I0(n5158), .I1(n5157), .I2(n4364), .I3(n5161), 
            .O(n5162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8774.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8775 (.I0(\i14/fifo_inst/buff[68][7] ), .I1(\i14/fifo_inst/buff[70][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8775.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8776 (.I0(\i14/fifo_inst/buff[71][7] ), .I1(\i14/fifo_inst/buff[69][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8776.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8777 (.I0(n5163), .I1(n5164), .I2(\fifo_inst/rd_index[3] ), 
            .I3(n4355), .O(n5165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8777.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8778 (.I0(n4358), .I1(n5156), .I2(n5165), .I3(n5162), 
            .O(n5166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__8778.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__8779 (.I0(\i14/fifo_inst/buff[84][7] ), .I1(\i14/fifo_inst/buff[86][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8779.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8780 (.I0(\i14/fifo_inst/buff[87][7] ), .I1(\i14/fifo_inst/buff[85][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8780.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8781 (.I0(\i14/fifo_inst/buff[80][7] ), .I1(\i14/fifo_inst/buff[82][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8781.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8782 (.I0(\i14/fifo_inst/buff[83][7] ), .I1(\i14/fifo_inst/buff[81][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n5169), .O(n5170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8782.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8783 (.I0(n5168), .I1(n5167), .I2(n5170), .I3(n4355), 
            .O(n5171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__8783.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__8784 (.I0(\i14/fifo_inst/buff[93][7] ), .I1(\i14/fifo_inst/buff[92][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcffa */ ;
    defparam LUT__8784.LUTMASK = 16'hcffa;
    EFX_LUT4 LUT__8785 (.I0(\i14/fifo_inst/buff[88][7] ), .I1(\i14/fifo_inst/buff[90][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__8785.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__8786 (.I0(\i14/fifo_inst/buff[91][7] ), .I1(\i14/fifo_inst/buff[89][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n5173), .O(n5174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__8786.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__8787 (.I0(\i14/fifo_inst/buff[94][7] ), .I1(\i14/fifo_inst/buff[95][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfacf */ ;
    defparam LUT__8787.LUTMASK = 16'hfacf;
    EFX_LUT4 LUT__8788 (.I0(n5172), .I1(n5175), .I2(n5174), .I3(n4355), 
            .O(n5176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__8788.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__8789 (.I0(n5176), .I1(n5171), .I2(n4475), .O(n5177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__8789.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__8790 (.I0(n5177), .I1(n5166), .I2(n4854), .I3(n4373), 
            .O(n5178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__8790.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__8791 (.I0(\i14/fifo_inst/buff[107][7] ), .I1(\i14/fifo_inst/buff[105][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8791.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8792 (.I0(\i14/fifo_inst/buff[104][7] ), .I1(\i14/fifo_inst/buff[106][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8792.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8793 (.I0(\i14/fifo_inst/buff[108][7] ), .I1(\i14/fifo_inst/buff[110][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8793.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8794 (.I0(\i14/fifo_inst/buff[111][7] ), .I1(\i14/fifo_inst/buff[109][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8794.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8795 (.I0(n5181), .I1(n5182), .I2(n4355), .O(n5183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8795.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8796 (.I0(n5180), .I1(n4355), .I2(n5179), .I3(n5183), 
            .O(n5184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8796.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8797 (.I0(\i14/fifo_inst/buff[99][7] ), .I1(\i14/fifo_inst/buff[97][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8797.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8798 (.I0(\i14/fifo_inst/buff[96][7] ), .I1(\i14/fifo_inst/buff[98][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8798.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8799 (.I0(\i14/fifo_inst/buff[100][7] ), .I1(\i14/fifo_inst/buff[102][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__8799.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__8800 (.I0(\i14/fifo_inst/buff[103][7] ), .I1(\i14/fifo_inst/buff[101][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(n5187), .O(n5188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__8800.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__8801 (.I0(n5186), .I1(n5185), .I2(n5188), .I3(n4355), 
            .O(n5189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__8801.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__8802 (.I0(n5189), .I1(n5184), .I2(n4373), .I3(n4475), 
            .O(n5190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8802.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8803 (.I0(\i14/fifo_inst/buff[123][7] ), .I1(\i14/fifo_inst/buff[121][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8803.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8804 (.I0(\i14/fifo_inst/buff[120][7] ), .I1(\i14/fifo_inst/buff[122][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8804.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8805 (.I0(\i14/fifo_inst/buff[127][7] ), .I1(\i14/fifo_inst/buff[125][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8805.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8806 (.I0(n5191), .I1(n5192), .I2(n5193), .I3(n4355), 
            .O(n5194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__8806.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__8807 (.I0(\i14/fifo_inst/buff[124][7] ), .I1(\i14/fifo_inst/buff[126][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8807.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8808 (.I0(n5195), .I1(n4355), .I2(n4475), .I3(n5194), 
            .O(n5196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0c */ ;
    defparam LUT__8808.LUTMASK = 16'h0b0c;
    EFX_LUT4 LUT__8809 (.I0(\i14/fifo_inst/buff[116][7] ), .I1(\i14/fifo_inst/buff[118][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8809.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8810 (.I0(\i14/fifo_inst/buff[119][7] ), .I1(\i14/fifo_inst/buff[117][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8810.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8811 (.I0(\i14/fifo_inst/buff[112][7] ), .I1(\i14/fifo_inst/buff[114][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8811.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8812 (.I0(\i14/fifo_inst/buff[115][7] ), .I1(\i14/fifo_inst/buff[113][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8812.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8813 (.I0(n5200), .I1(n4355), .I2(n5199), .I3(n4475), 
            .O(n5201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8813.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8814 (.I0(n5197), .I1(n5198), .I2(n4355), .I3(n5201), 
            .O(n5202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8814.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8815 (.I0(n5196), .I1(n5202), .I2(n4373), .I3(n4888), 
            .O(n5203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8815.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8816 (.I0(\i14/fifo_inst/buff[52][7] ), .I1(\i14/fifo_inst/buff[54][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8816.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8817 (.I0(\i14/fifo_inst/buff[55][7] ), .I1(\i14/fifo_inst/buff[53][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8817.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8818 (.I0(\i14/fifo_inst/buff[51][7] ), .I1(\i14/fifo_inst/buff[49][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8818.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8819 (.I0(\i14/fifo_inst/buff[48][7] ), .I1(\i14/fifo_inst/buff[50][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8819.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8820 (.I0(n5207), .I1(n4355), .I2(n5206), .I3(n4475), 
            .O(n5208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8820.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8821 (.I0(n5204), .I1(n5205), .I2(n4355), .I3(n5208), 
            .O(n5209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8821.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8822 (.I0(\i14/fifo_inst/buff[59][7] ), .I1(\i14/fifo_inst/buff[57][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8822.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8823 (.I0(\i14/fifo_inst/buff[56][7] ), .I1(\i14/fifo_inst/buff[58][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8823.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8824 (.I0(\i14/fifo_inst/buff[60][7] ), .I1(\i14/fifo_inst/buff[62][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8824.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8825 (.I0(\i14/fifo_inst/buff[63][7] ), .I1(\i14/fifo_inst/buff[61][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8825.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8826 (.I0(n5212), .I1(n5213), .I2(n4355), .I3(n4475), 
            .O(n5214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8826.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8827 (.I0(n5211), .I1(n4355), .I2(n5210), .I3(n5214), 
            .O(n5215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8827.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8828 (.I0(n5209), .I1(n5215), .I2(n4373), .O(n5216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8828.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8829 (.I0(\i14/fifo_inst/buff[32][7] ), .I1(\i14/fifo_inst/buff[34][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8829.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8830 (.I0(\i14/fifo_inst/buff[35][7] ), .I1(\i14/fifo_inst/buff[33][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8830.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8831 (.I0(\i14/fifo_inst/buff[36][7] ), .I1(\i14/fifo_inst/buff[38][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8831.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8832 (.I0(\i14/fifo_inst/buff[39][7] ), .I1(\i14/fifo_inst/buff[37][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8832.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8833 (.I0(n5219), .I1(n5220), .I2(n4355), .I3(n4475), 
            .O(n5221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__8833.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__8834 (.I0(n5218), .I1(n4355), .I2(n5217), .I3(n5221), 
            .O(n5222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8834.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8835 (.I0(\i14/fifo_inst/buff[40][7] ), .I1(\i14/fifo_inst/buff[42][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8835.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8836 (.I0(\i14/fifo_inst/buff[43][7] ), .I1(\i14/fifo_inst/buff[41][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8836.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8837 (.I0(\i14/fifo_inst/buff[44][7] ), .I1(\i14/fifo_inst/buff[46][7] ), 
            .I2(\fifo_inst/rd_index[1] ), .I3(\fifo_inst/rd_index[0] ), 
            .O(n5225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8837.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8838 (.I0(\i14/fifo_inst/buff[47][7] ), .I1(\i14/fifo_inst/buff[45][7] ), 
            .I2(\fifo_inst/rd_index[0] ), .I3(\fifo_inst/rd_index[1] ), 
            .O(n5226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8838.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8839 (.I0(n5225), .I1(n5226), .I2(n4355), .I3(n4475), 
            .O(n5227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8839.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8840 (.I0(n5224), .I1(n4355), .I2(n5223), .I3(n5227), 
            .O(n5228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8840.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8841 (.I0(n5228), .I1(n4373), .I2(n5222), .I3(n4913), 
            .O(n5229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8841.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8842 (.I0(n5216), .I1(n5229), .I2(n5190), .I3(n5203), 
            .O(n5230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__8842.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__8843 (.I0(n4809), .I1(\rx_d[7] ), .O(n5231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8843.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8844 (.I0(n5178), .I1(n5154), .I2(n5230), .I3(n5231), 
            .O(\fifo_inst/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10 */ ;
    defparam LUT__8844.LUTMASK = 16'hff10;
    EFX_LUT4 LUT__8845 (.I0(\reg_addr[2] ), .I1(n4318), .I2(n4239), .I3(\reg_addr[1] ), 
            .O(rx_en_tx_packet_len)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__8845.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__8846 (.I0(rx_en_tx_packet_len), .I1(\tx_fifo/wr_index[0] ), 
            .O(\tx_fifo/n153 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8846.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8847 (.I0(\tx_fifo/sync_wr[1] ), .I1(\tx_fifo/sync_wr[0] ), 
            .O(n5232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8847.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8848 (.I0(rx_en_tx_packet_len), .I1(n5232), .O(ceg_net234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8848.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8849 (.I0(rx_en_tx_packet_len), .I1(\tx_fifo/rd_index[0] ), 
            .O(\tx_fifo/n162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8849.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8850 (.I0(n5232), .I1(\tx_fifo/sync_rd[0] ), .I2(\tx_fifo/sync_rd[1] ), 
            .O(n5233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8850.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8851 (.I0(\tx_fifo/wr_index[6] ), .I1(\tx_fifo/rd_index[6] ), 
            .I2(\tx_fifo/wr_index[7] ), .I3(\tx_fifo/rd_index[7] ), .O(n5234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__8851.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__8852 (.I0(\tx_fifo/wr_index[2] ), .I1(\tx_fifo/rd_index[2] ), 
            .I2(\tx_fifo/wr_index[3] ), .I3(\tx_fifo/rd_index[3] ), .O(n5235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__8852.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__8853 (.I0(\tx_fifo/wr_index[0] ), .I1(\tx_fifo/rd_index[0] ), 
            .I2(\tx_fifo/wr_index[1] ), .I3(\tx_fifo/rd_index[1] ), .O(n5236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__8853.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__8854 (.I0(\tx_fifo/wr_index[4] ), .I1(\tx_fifo/rd_index[4] ), 
            .I2(\tx_fifo/wr_index[5] ), .I3(\tx_fifo/rd_index[5] ), .O(n5237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__8854.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__8855 (.I0(n5234), .I1(n5235), .I2(n5236), .I3(n5237), 
            .O(n5238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8855.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8856 (.I0(n5238), .I1(n5233), .I2(rx_en_tx_packet_len), 
            .O(ceg_net252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__8856.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__8857 (.I0(rx_en_tx_packet_len), .I1(\rx_d[0] ), .O(\data_to_tx_packet_len_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8857.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8858 (.I0(\reg_addr[2] ), .I1(n4343), .I2(n4239), .I3(\reg_addr[1] ), 
            .O(rx_en_tx_packet)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__8858.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__8859 (.I0(n4245), .I1(\reg_addr[0] ), .O(tx_en_tx_packet)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8859.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8860 (.I0(\i15/tx_fifo/buff[75][0] ), .I1(\i15/tx_fifo/buff[73][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8860.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8861 (.I0(\i15/tx_fifo/buff[72][0] ), .I1(\i15/tx_fifo/buff[74][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8861.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8862 (.I0(\tx_fifo/rd_index[0] ), .I1(\tx_fifo/rd_index[1] ), 
            .I2(\tx_fifo/rd_index[2] ), .O(n5241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__8862.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__8863 (.I0(\i15/tx_fifo/buff[76][0] ), .I1(\i15/tx_fifo/buff[78][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8863.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8864 (.I0(\i15/tx_fifo/buff[79][0] ), .I1(\i15/tx_fifo/buff[77][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__8864.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__8865 (.I0(n5243), .I1(n5242), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__8865.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__8866 (.I0(n5240), .I1(n5241), .I2(n5239), .I3(n5244), 
            .O(n5245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8866.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8867 (.I0(\i15/tx_fifo/buff[67][0] ), .I1(\i15/tx_fifo/buff[65][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8867.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8868 (.I0(\i15/tx_fifo/buff[64][0] ), .I1(\i15/tx_fifo/buff[66][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8868.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8869 (.I0(\i15/tx_fifo/buff[68][0] ), .I1(\i15/tx_fifo/buff[70][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8869.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8870 (.I0(\i15/tx_fifo/buff[71][0] ), .I1(\i15/tx_fifo/buff[69][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__8870.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__8871 (.I0(n5249), .I1(n5248), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__8871.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__8872 (.I0(n5247), .I1(n5241), .I2(n5246), .I3(n5250), 
            .O(n5251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8872.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8873 (.I0(\tx_fifo/rd_index[0] ), .I1(\tx_fifo/rd_index[1] ), 
            .I2(\tx_fifo/rd_index[2] ), .I3(\tx_fifo/rd_index[3] ), .O(n5252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h807f */ ;
    defparam LUT__8873.LUTMASK = 16'h807f;
    EFX_LUT4 LUT__8874 (.I0(n5251), .I1(n5245), .I2(n5252), .O(n5253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8874.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8875 (.I0(\i15/tx_fifo/buff[83][0] ), .I1(\i15/tx_fifo/buff[81][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8875.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8876 (.I0(\i15/tx_fifo/buff[80][0] ), .I1(\i15/tx_fifo/buff[82][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8876.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8877 (.I0(\i15/tx_fifo/buff[84][0] ), .I1(\i15/tx_fifo/buff[86][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8877.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8878 (.I0(\i15/tx_fifo/buff[87][0] ), .I1(\i15/tx_fifo/buff[85][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8878.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8879 (.I0(n5257), .I1(n5256), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__8879.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__8880 (.I0(n5255), .I1(n5241), .I2(n5254), .I3(n5258), 
            .O(n5259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8880.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8881 (.I0(\i15/tx_fifo/buff[91][0] ), .I1(\i15/tx_fifo/buff[89][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8881.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8882 (.I0(\i15/tx_fifo/buff[88][0] ), .I1(\i15/tx_fifo/buff[90][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8882.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8883 (.I0(\i15/tx_fifo/buff[92][0] ), .I1(\i15/tx_fifo/buff[94][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8883.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8884 (.I0(\i15/tx_fifo/buff[95][0] ), .I1(\i15/tx_fifo/buff[93][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__8884.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__8885 (.I0(n5263), .I1(n5262), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__8885.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__8886 (.I0(n5261), .I1(n5241), .I2(n5260), .I3(n5264), 
            .O(n5265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8886.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8887 (.I0(n5265), .I1(n5259), .I2(n5252), .O(n5266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__8887.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__8888 (.I0(\tx_fifo/rd_index[0] ), .I1(\tx_fifo/rd_index[1] ), 
            .I2(\tx_fifo/rd_index[2] ), .I3(\tx_fifo/rd_index[3] ), .O(n5267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__8888.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__8889 (.I0(n5267), .I1(\tx_fifo/rd_index[4] ), .O(n5268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8889.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8890 (.I0(n5268), .I1(\tx_fifo/rd_index[5] ), .I2(\tx_fifo/rd_index[6] ), 
            .O(n5269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7e7 */ ;
    defparam LUT__8890.LUTMASK = 16'he7e7;
    EFX_LUT4 LUT__8891 (.I0(n5267), .I1(\tx_fifo/rd_index[4] ), .O(n5270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__8891.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__8892 (.I0(n5266), .I1(n5253), .I2(n5269), .I3(n5270), 
            .O(n5271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8892.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8893 (.I0(\i15/tx_fifo/buff[47][0] ), .I1(\i15/tx_fifo/buff[45][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8893.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8894 (.I0(\i15/tx_fifo/buff[44][0] ), .I1(\i15/tx_fifo/buff[46][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8894.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8895 (.I0(n5272), .I1(n5273), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__8895.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__8896 (.I0(\i15/tx_fifo/buff[40][0] ), .I1(\i15/tx_fifo/buff[42][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8896.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8897 (.I0(\i15/tx_fifo/buff[43][0] ), .I1(\i15/tx_fifo/buff[41][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8897.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8898 (.I0(\tx_fifo/rd_index[0] ), .I1(\tx_fifo/rd_index[1] ), 
            .I2(\tx_fifo/rd_index[3] ), .I3(\tx_fifo/rd_index[2] ), .O(n5277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf78f */ ;
    defparam LUT__8898.LUTMASK = 16'hf78f;
    EFX_LUT4 LUT__8899 (.I0(n5276), .I1(n5275), .I2(n5277), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8899.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8900 (.I0(\i15/tx_fifo/buff[32][0] ), .I1(\i15/tx_fifo/buff[34][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8900.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8901 (.I0(\i15/tx_fifo/buff[35][0] ), .I1(\i15/tx_fifo/buff[33][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8901.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8902 (.I0(\tx_fifo/rd_index[0] ), .I1(\tx_fifo/rd_index[1] ), 
            .I2(\tx_fifo/rd_index[2] ), .I3(\tx_fifo/rd_index[3] ), .O(n5281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ff8 */ ;
    defparam LUT__8902.LUTMASK = 16'h7ff8;
    EFX_LUT4 LUT__8903 (.I0(n5280), .I1(n5279), .I2(n5281), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8903.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8904 (.I0(\i15/tx_fifo/buff[36][0] ), .I1(\i15/tx_fifo/buff[38][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8904.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8905 (.I0(\i15/tx_fifo/buff[39][0] ), .I1(\i15/tx_fifo/buff[37][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8905.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8906 (.I0(n5283), .I1(n5284), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8906.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8907 (.I0(n5274), .I1(n5278), .I2(n5282), .I3(n5285), 
            .O(n5286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8907.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8908 (.I0(\i15/tx_fifo/buff[55][0] ), .I1(\i15/tx_fifo/buff[53][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8908.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8909 (.I0(\i15/tx_fifo/buff[52][0] ), .I1(\i15/tx_fifo/buff[54][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8909.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8910 (.I0(\i15/tx_fifo/buff[48][0] ), .I1(\i15/tx_fifo/buff[50][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8910.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8911 (.I0(\i15/tx_fifo/buff[51][0] ), .I1(\i15/tx_fifo/buff[49][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__8911.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__8912 (.I0(n5290), .I1(n5289), .I2(n5241), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__8912.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__8913 (.I0(n5287), .I1(n5288), .I2(n5241), .I3(n5291), 
            .O(n5292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8913.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8914 (.I0(\i15/tx_fifo/buff[63][0] ), .I1(\i15/tx_fifo/buff[61][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8914.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8915 (.I0(\i15/tx_fifo/buff[60][0] ), .I1(\i15/tx_fifo/buff[62][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8915.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8916 (.I0(\i15/tx_fifo/buff[56][0] ), .I1(\i15/tx_fifo/buff[58][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8916.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8917 (.I0(\i15/tx_fifo/buff[59][0] ), .I1(\i15/tx_fifo/buff[57][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8917.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8918 (.I0(n5296), .I1(n5295), .I2(n5241), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__8918.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__8919 (.I0(n5293), .I1(n5294), .I2(n5241), .I3(n5297), 
            .O(n5298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__8919.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__8920 (.I0(n5298), .I1(n5292), .I2(n5252), .O(n5299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__8920.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__8921 (.I0(\tx_fifo/rd_index[6] ), .I1(n5268), .I2(\tx_fifo/rd_index[5] ), 
            .O(n5300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__8921.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__8922 (.I0(n5299), .I1(n5286), .I2(n5270), .I3(n5300), 
            .O(n5301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__8922.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__8923 (.I0(n5268), .I1(\tx_fifo/rd_index[5] ), .I2(\tx_fifo/rd_index[6] ), 
            .O(n5302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__8923.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__8924 (.I0(n5270), .I1(n5302), .O(n5303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8924.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8925 (.I0(\i15/tx_fifo/buff[99][0] ), .I1(\i15/tx_fifo/buff[97][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8925.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8926 (.I0(\i15/tx_fifo/buff[96][0] ), .I1(\i15/tx_fifo/buff[98][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8926.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8927 (.I0(\i15/tx_fifo/buff[100][0] ), .I1(\i15/tx_fifo/buff[102][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8927.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8928 (.I0(\i15/tx_fifo/buff[103][0] ), .I1(\i15/tx_fifo/buff[101][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__8928.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__8929 (.I0(n5307), .I1(n5306), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__8929.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__8930 (.I0(n5305), .I1(n5241), .I2(n5304), .I3(n5308), 
            .O(n5309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8930.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8931 (.I0(\i15/tx_fifo/buff[107][0] ), .I1(\i15/tx_fifo/buff[105][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8931.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8932 (.I0(\i15/tx_fifo/buff[104][0] ), .I1(\i15/tx_fifo/buff[106][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8932.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8933 (.I0(\i15/tx_fifo/buff[108][0] ), .I1(\i15/tx_fifo/buff[110][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8933.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8934 (.I0(\i15/tx_fifo/buff[111][0] ), .I1(\i15/tx_fifo/buff[109][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__8934.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__8935 (.I0(n5313), .I1(n5312), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__8935.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__8936 (.I0(n5311), .I1(n5241), .I2(n5310), .I3(n5314), 
            .O(n5315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8936.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8937 (.I0(n5315), .I1(n5309), .I2(n5252), .O(n5316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__8937.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__8938 (.I0(\i15/tx_fifo/buff[23][0] ), .I1(\i15/tx_fifo/buff[21][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8938.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8939 (.I0(\i15/tx_fifo/buff[20][0] ), .I1(\i15/tx_fifo/buff[22][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8939.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8940 (.I0(n5317), .I1(n5318), .I2(n5241), .O(n5319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8940.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8941 (.I0(\i15/tx_fifo/buff[19][0] ), .I1(\i15/tx_fifo/buff[17][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8941.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8942 (.I0(\i15/tx_fifo/buff[16][0] ), .I1(\i15/tx_fifo/buff[18][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8942.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8943 (.I0(n5321), .I1(n5241), .I2(n5320), .I3(n5252), 
            .O(n5322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__8943.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__8944 (.I0(\i15/tx_fifo/buff[31][0] ), .I1(\i15/tx_fifo/buff[29][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8944.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8945 (.I0(\i15/tx_fifo/buff[28][0] ), .I1(\i15/tx_fifo/buff[30][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8945.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8946 (.I0(n5323), .I1(n5324), .I2(n5241), .O(n5325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8946.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8947 (.I0(\i15/tx_fifo/buff[27][0] ), .I1(\i15/tx_fifo/buff[25][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8947.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8948 (.I0(\i15/tx_fifo/buff[24][0] ), .I1(\i15/tx_fifo/buff[26][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8948.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8949 (.I0(n5327), .I1(n5241), .I2(n5326), .I3(n5252), 
            .O(n5328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__8949.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__8950 (.I0(n5325), .I1(n5328), .I2(n5319), .I3(n5322), 
            .O(n5329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__8950.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__8951 (.I0(n5267), .I1(\tx_fifo/rd_index[4] ), .I2(\tx_fifo/rd_index[5] ), 
            .I3(\tx_fifo/rd_index[6] ), .O(n5330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ff8 */ ;
    defparam LUT__8951.LUTMASK = 16'h7ff8;
    EFX_LUT4 LUT__8952 (.I0(n5330), .I1(n5270), .O(n5331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8952.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8953 (.I0(\i15/tx_fifo/buff[11][0] ), .I1(\i15/tx_fifo/buff[9][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8953.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8954 (.I0(\i15/tx_fifo/buff[8][0] ), .I1(\i15/tx_fifo/buff[10][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8954.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8955 (.I0(\i15/tx_fifo/buff[12][0] ), .I1(\i15/tx_fifo/buff[14][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8955.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8956 (.I0(n5332), .I1(n5333), .I2(n5334), .I3(n5241), 
            .O(n5335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__8956.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__8957 (.I0(\i15/tx_fifo/buff[15][0] ), .I1(\i15/tx_fifo/buff[13][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8957.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8958 (.I0(n5336), .I1(n5241), .I2(n5335), .I3(n5252), 
            .O(n5337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__8958.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__8959 (.I0(\i15/tx_fifo/buff[7][0] ), .I1(\i15/tx_fifo/buff[5][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8959.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8960 (.I0(\i15/tx_fifo/buff[4][0] ), .I1(\i15/tx_fifo/buff[6][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8960.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8961 (.I0(n5338), .I1(n5339), .I2(n5241), .O(n5340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__8961.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__8962 (.I0(\i15/tx_fifo/buff[3][0] ), .I1(\i15/tx_fifo/buff[1][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8962.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8963 (.I0(\i15/tx_fifo/buff[0][0] ), .I1(\i15/tx_fifo/buff[2][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8963.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8964 (.I0(n5341), .I1(n5342), .I2(n5241), .O(n5343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8964.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8965 (.I0(n5267), .I1(\tx_fifo/rd_index[4] ), .I2(\tx_fifo/rd_index[5] ), 
            .I3(\tx_fifo/rd_index[6] ), .O(n5344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ffe */ ;
    defparam LUT__8965.LUTMASK = 16'h7ffe;
    EFX_LUT4 LUT__8966 (.I0(n5343), .I1(n5340), .I2(n5252), .I3(n5344), 
            .O(n5345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__8966.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__8967 (.I0(n5337), .I1(n5345), .I2(n5329), .I3(n5331), 
            .O(n5346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__8967.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__8968 (.I0(\i15/tx_fifo/buff[112][0] ), .I1(\i15/tx_fifo/buff[114][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__8968.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__8969 (.I0(\i15/tx_fifo/buff[115][0] ), .I1(\i15/tx_fifo/buff[113][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__8969.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__8970 (.I0(n5348), .I1(n5347), .I2(n5281), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__8970.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__8971 (.I0(\i15/tx_fifo/buff[119][0] ), .I1(\i15/tx_fifo/buff[117][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8971.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8972 (.I0(\i15/tx_fifo/buff[116][0] ), .I1(\i15/tx_fifo/buff[118][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8972.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8973 (.I0(n5350), .I1(n5351), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__8973.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__8974 (.I0(\i15/tx_fifo/buff[127][0] ), .I1(\i15/tx_fifo/buff[125][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8974.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8975 (.I0(\i15/tx_fifo/buff[124][0] ), .I1(\i15/tx_fifo/buff[126][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8975.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8976 (.I0(n5353), .I1(n5354), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__8976.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__8977 (.I0(\i15/tx_fifo/buff[123][0] ), .I1(\i15/tx_fifo/buff[121][0] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__8977.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__8978 (.I0(\i15/tx_fifo/buff[120][0] ), .I1(\i15/tx_fifo/buff[122][0] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__8978.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__8979 (.I0(n5277), .I1(n5356), .I2(n5357), .O(n5358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8979.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8980 (.I0(n5349), .I1(n5352), .I2(n5355), .I3(n5358), 
            .O(n5359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__8980.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__8981 (.I0(n5270), .I1(\tx_fifo/rd_index[5] ), .I2(\tx_fifo/rd_index[6] ), 
            .O(n5360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__8981.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__8982 (.I0(rx_en_tx_packet_len), .I1(n5238), .I2(n5232), 
            .O(n5361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__8982.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__8983 (.I0(n5360), .I1(n5359), .I2(n5361), .O(n5362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__8983.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__8984 (.I0(n5316), .I1(n5303), .I2(n5346), .I3(n5362), 
            .O(n5363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__8984.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__8985 (.I0(rx_en_tx_packet), .I1(\rx_d[0] ), .O(\data_to_tx_packet_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8985.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8986 (.I0(\data_to_tx_packet_reg[0] ), .I1(n5232), .O(n5364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__8986.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__8987 (.I0(n5301), .I1(n5271), .I2(n5363), .I3(n5364), 
            .O(\tx_fifo/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10 */ ;
    defparam LUT__8987.LUTMASK = 16'hff10;
    EFX_LUT4 LUT__8988 (.I0(n5238), .I1(n5232), .I2(n5233), .I3(rx_en_tx_packet_len), 
            .O(ceg_net458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__8988.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__8989 (.I0(rx_en_tx_packet_len), .I1(n147), .O(\tx_fifo/n152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8989.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8990 (.I0(rx_en_tx_packet_len), .I1(n3219), .O(\tx_fifo/n151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8990.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8991 (.I0(rx_en_tx_packet_len), .I1(n3215), .O(\tx_fifo/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8991.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8992 (.I0(rx_en_tx_packet_len), .I1(n3212), .O(\tx_fifo/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8992.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8993 (.I0(rx_en_tx_packet_len), .I1(n3208), .O(\tx_fifo/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8993.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8994 (.I0(rx_en_tx_packet_len), .I1(n3205), .O(\tx_fifo/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8994.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8995 (.I0(rx_en_tx_packet_len), .I1(n3202), .O(\tx_fifo/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8995.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8996 (.I0(rx_en_tx_packet_len), .I1(\tx_fifo/rd_index[0] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(\tx_fifo/n161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__8996.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__8997 (.I0(rx_en_tx_packet_len), .I1(n5241), .O(\tx_fifo/n160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8997.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__8998 (.I0(rx_en_tx_packet_len), .I1(n5252), .O(\tx_fifo/n159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__8998.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__8999 (.I0(rx_en_tx_packet_len), .I1(n5270), .O(\tx_fifo/n158 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__8999.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9000 (.I0(rx_en_tx_packet_len), .I1(n5268), .I2(\tx_fifo/rd_index[5] ), 
            .O(\tx_fifo/n157 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__9000.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__9001 (.I0(n5268), .I1(\tx_fifo/rd_index[5] ), .I2(rx_en_tx_packet_len), 
            .I3(\tx_fifo/rd_index[6] ), .O(\tx_fifo/n156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__9001.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__9002 (.I0(n5268), .I1(\tx_fifo/rd_index[5] ), .I2(\tx_fifo/rd_index[6] ), 
            .I3(\tx_fifo/rd_index[7] ), .O(n5365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h807f */ ;
    defparam LUT__9002.LUTMASK = 16'h807f;
    EFX_LUT4 LUT__9003 (.I0(rx_en_tx_packet_len), .I1(n5365), .O(\tx_fifo/n155 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__9003.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__9004 (.I0(rx_en_tx_packet_len), .I1(\rx_d[1] ), .O(\data_to_tx_packet_len_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9004.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9005 (.I0(rx_en_tx_packet_len), .I1(\rx_d[2] ), .O(\data_to_tx_packet_len_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9005.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9006 (.I0(rx_en_tx_packet_len), .I1(\rx_d[3] ), .O(\data_to_tx_packet_len_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9006.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9007 (.I0(rx_en_tx_packet_len), .I1(\rx_d[4] ), .O(\data_to_tx_packet_len_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9007.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9008 (.I0(rx_en_tx_packet_len), .I1(\rx_d[5] ), .O(\data_to_tx_packet_len_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9008.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9009 (.I0(rx_en_tx_packet_len), .I1(\rx_d[6] ), .O(\data_to_tx_packet_len_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9009.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9010 (.I0(rx_en_tx_packet_len), .I1(\rx_d[7] ), .O(\data_to_tx_packet_len_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9010.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9011 (.I0(\i15/tx_fifo/buff[4][1] ), .I1(\i15/tx_fifo/buff[6][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9011.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9012 (.I0(\i15/tx_fifo/buff[7][1] ), .I1(\i15/tx_fifo/buff[5][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9012.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9013 (.I0(n5367), .I1(n5366), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9013.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9014 (.I0(\i15/tx_fifo/buff[0][1] ), .I1(\i15/tx_fifo/buff[2][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9014.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9015 (.I0(\i15/tx_fifo/buff[3][1] ), .I1(\i15/tx_fifo/buff[1][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9015.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9016 (.I0(n5370), .I1(n5369), .I2(n5241), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9016.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9017 (.I0(\i15/tx_fifo/buff[15][1] ), .I1(\i15/tx_fifo/buff[13][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9017.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9018 (.I0(\i15/tx_fifo/buff[12][1] ), .I1(\i15/tx_fifo/buff[14][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9018.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9019 (.I0(\i15/tx_fifo/buff[11][1] ), .I1(\i15/tx_fifo/buff[9][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9019.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9020 (.I0(\i15/tx_fifo/buff[8][1] ), .I1(\i15/tx_fifo/buff[10][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9020.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9021 (.I0(n5375), .I1(n5241), .I2(n5374), .I3(n5252), 
            .O(n5376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9021.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9022 (.I0(n5372), .I1(n5373), .I2(n5241), .I3(n5376), 
            .O(n5377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9022.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9023 (.I0(n5371), .I1(n5368), .I2(n5252), .I3(n5377), 
            .O(n5378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9023.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9024 (.I0(\i15/tx_fifo/buff[24][1] ), .I1(\i15/tx_fifo/buff[26][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9024.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9025 (.I0(\i15/tx_fifo/buff[27][1] ), .I1(\i15/tx_fifo/buff[25][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5379), .O(n5380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9025.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9026 (.I0(\i15/tx_fifo/buff[31][1] ), .I1(\i15/tx_fifo/buff[29][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9026.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9027 (.I0(\i15/tx_fifo/buff[28][1] ), .I1(\i15/tx_fifo/buff[30][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9027.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9028 (.I0(n5381), .I1(n5382), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9028.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9029 (.I0(\i15/tx_fifo/buff[16][1] ), .I1(\i15/tx_fifo/buff[18][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9029.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9030 (.I0(\i15/tx_fifo/buff[19][1] ), .I1(\i15/tx_fifo/buff[17][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9030.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9031 (.I0(n5385), .I1(n5384), .I2(n5281), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9031.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9032 (.I0(\i15/tx_fifo/buff[23][1] ), .I1(\i15/tx_fifo/buff[21][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9032.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9033 (.I0(\i15/tx_fifo/buff[20][1] ), .I1(\i15/tx_fifo/buff[22][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9033.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9034 (.I0(n5387), .I1(n5388), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9034.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9035 (.I0(n5383), .I1(n5386), .I2(n5389), .I3(n5270), 
            .O(n5390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9035.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9036 (.I0(n5277), .I1(n5380), .I2(n5390), .I3(n5330), 
            .O(n5391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__9036.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__9037 (.I0(\i15/tx_fifo/buff[95][1] ), .I1(\i15/tx_fifo/buff[93][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9037.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9038 (.I0(\i15/tx_fifo/buff[92][1] ), .I1(\i15/tx_fifo/buff[94][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9038.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9039 (.I0(n5392), .I1(n5393), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9039.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9040 (.I0(\i15/tx_fifo/buff[83][1] ), .I1(\i15/tx_fifo/buff[81][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9040.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9041 (.I0(\i15/tx_fifo/buff[80][1] ), .I1(\i15/tx_fifo/buff[82][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9041.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9042 (.I0(n5281), .I1(n5395), .I2(n5396), .O(n5397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9042.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9043 (.I0(\i15/tx_fifo/buff[91][1] ), .I1(\i15/tx_fifo/buff[89][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9043.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9044 (.I0(\i15/tx_fifo/buff[88][1] ), .I1(\i15/tx_fifo/buff[90][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9044.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9045 (.I0(n5277), .I1(n5398), .I2(n5399), .O(n5400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9045.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9046 (.I0(\i15/tx_fifo/buff[87][1] ), .I1(\i15/tx_fifo/buff[85][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9046.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9047 (.I0(\i15/tx_fifo/buff[84][1] ), .I1(\i15/tx_fifo/buff[86][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9047.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9048 (.I0(n5401), .I1(n5402), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9048.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9049 (.I0(n5394), .I1(n5397), .I2(n5400), .I3(n5403), 
            .O(n5404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9049.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9050 (.I0(\i15/tx_fifo/buff[71][1] ), .I1(\i15/tx_fifo/buff[69][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9050.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9051 (.I0(\i15/tx_fifo/buff[68][1] ), .I1(\i15/tx_fifo/buff[70][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9051.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9052 (.I0(n5405), .I1(n5406), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9052.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9053 (.I0(\i15/tx_fifo/buff[67][1] ), .I1(\i15/tx_fifo/buff[65][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9053.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9054 (.I0(\i15/tx_fifo/buff[64][1] ), .I1(\i15/tx_fifo/buff[66][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9054.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9055 (.I0(n5281), .I1(n5408), .I2(n5409), .O(n5410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9055.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9056 (.I0(\i15/tx_fifo/buff[75][1] ), .I1(\i15/tx_fifo/buff[73][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9056.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9057 (.I0(\i15/tx_fifo/buff[72][1] ), .I1(\i15/tx_fifo/buff[74][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9057.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9058 (.I0(n5277), .I1(n5411), .I2(n5412), .O(n5413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9058.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9059 (.I0(\i15/tx_fifo/buff[79][1] ), .I1(\i15/tx_fifo/buff[77][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9059.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9060 (.I0(\i15/tx_fifo/buff[76][1] ), .I1(\i15/tx_fifo/buff[78][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9060.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9061 (.I0(n5414), .I1(n5415), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9061.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9062 (.I0(n5407), .I1(n5410), .I2(n5413), .I3(n5416), 
            .O(n5417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9062.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9063 (.I0(n5417), .I1(n5404), .I2(n5269), .I3(n5270), 
            .O(n5418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__9063.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__9064 (.I0(n5270), .I1(n5378), .I2(n5391), .I3(n5418), 
            .O(n5419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__9064.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__9065 (.I0(\i15/tx_fifo/buff[123][1] ), .I1(\i15/tx_fifo/buff[121][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9065.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9066 (.I0(\i15/tx_fifo/buff[120][1] ), .I1(\i15/tx_fifo/buff[122][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9066.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9067 (.I0(\i15/tx_fifo/buff[127][1] ), .I1(\i15/tx_fifo/buff[125][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9067.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9068 (.I0(\i15/tx_fifo/buff[124][1] ), .I1(\i15/tx_fifo/buff[126][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9068.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9069 (.I0(n5422), .I1(n5423), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9069.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9070 (.I0(\i15/tx_fifo/buff[119][1] ), .I1(\i15/tx_fifo/buff[117][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9070.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9071 (.I0(\i15/tx_fifo/buff[116][1] ), .I1(\i15/tx_fifo/buff[118][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9071.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9072 (.I0(n5425), .I1(n5426), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9072.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9073 (.I0(\i15/tx_fifo/buff[115][1] ), .I1(\i15/tx_fifo/buff[113][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9073.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9074 (.I0(\i15/tx_fifo/buff[112][1] ), .I1(\i15/tx_fifo/buff[114][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9074.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9075 (.I0(n5281), .I1(n5428), .I2(n5429), .O(n5430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9075.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9076 (.I0(n5424), .I1(n5427), .I2(n5430), .I3(n5270), 
            .O(n5431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9076.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9077 (.I0(n5420), .I1(n5421), .I2(n5277), .I3(n5431), 
            .O(n5432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9077.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9078 (.I0(\i15/tx_fifo/buff[111][1] ), .I1(\i15/tx_fifo/buff[109][1] ), 
            .I2(\tx_fifo/rd_index[3] ), .I3(\tx_fifo/rd_index[1] ), .O(n5433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__9078.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__9079 (.I0(\i15/tx_fifo/buff[103][1] ), .I1(\i15/tx_fifo/buff[101][1] ), 
            .I2(\tx_fifo/rd_index[3] ), .I3(n5433), .O(n5434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__9079.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__9080 (.I0(\i15/tx_fifo/buff[100][1] ), .I1(\i15/tx_fifo/buff[102][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9080.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9081 (.I0(\i15/tx_fifo/buff[108][1] ), .I1(\i15/tx_fifo/buff[110][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9081.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9082 (.I0(n5435), .I1(n5436), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__9082.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__9083 (.I0(\i15/tx_fifo/buff[96][1] ), .I1(\i15/tx_fifo/buff[98][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9083.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9084 (.I0(\i15/tx_fifo/buff[99][1] ), .I1(\i15/tx_fifo/buff[97][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5438), .O(n5439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9084.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9085 (.I0(\i15/tx_fifo/buff[107][1] ), .I1(\i15/tx_fifo/buff[105][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9085.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9086 (.I0(\i15/tx_fifo/buff[104][1] ), .I1(\i15/tx_fifo/buff[106][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9086.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9087 (.I0(n5277), .I1(n5440), .I2(n5441), .O(n5442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9087.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9088 (.I0(n5281), .I1(n5439), .I2(n5270), .I3(n5442), 
            .O(n5443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__9088.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__9089 (.I0(n5434), .I1(\tx_fifo/rd_index[0] ), .I2(n5437), 
            .I3(n5443), .O(n5444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__9089.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__9090 (.I0(\i15/tx_fifo/buff[63][1] ), .I1(\i15/tx_fifo/buff[61][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9090.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9091 (.I0(\i15/tx_fifo/buff[60][1] ), .I1(\i15/tx_fifo/buff[62][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9091.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9092 (.I0(n5445), .I1(n5446), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9092.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9093 (.I0(\i15/tx_fifo/buff[55][1] ), .I1(\i15/tx_fifo/buff[53][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9093.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9094 (.I0(\i15/tx_fifo/buff[52][1] ), .I1(\i15/tx_fifo/buff[54][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9094.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9095 (.I0(n5448), .I1(n5449), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9095.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9096 (.I0(\i15/tx_fifo/buff[59][1] ), .I1(\i15/tx_fifo/buff[57][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9096.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9097 (.I0(\i15/tx_fifo/buff[56][1] ), .I1(\i15/tx_fifo/buff[58][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9097.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9098 (.I0(n5277), .I1(n5451), .I2(n5452), .O(n5453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9098.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9099 (.I0(\i15/tx_fifo/buff[51][1] ), .I1(\i15/tx_fifo/buff[49][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9099.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9100 (.I0(\i15/tx_fifo/buff[48][1] ), .I1(\i15/tx_fifo/buff[50][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9100.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9101 (.I0(n5281), .I1(n5454), .I2(n5455), .O(n5456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9101.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9102 (.I0(n5447), .I1(n5450), .I2(n5453), .I3(n5456), 
            .O(n5457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9102.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9103 (.I0(\i15/tx_fifo/buff[39][1] ), .I1(\i15/tx_fifo/buff[37][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9103.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9104 (.I0(\i15/tx_fifo/buff[36][1] ), .I1(\i15/tx_fifo/buff[38][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9104.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9105 (.I0(n5458), .I1(n5459), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9105.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9106 (.I0(\i15/tx_fifo/buff[47][1] ), .I1(\i15/tx_fifo/buff[45][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9106.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9107 (.I0(\i15/tx_fifo/buff[44][1] ), .I1(\i15/tx_fifo/buff[46][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9107.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9108 (.I0(n5461), .I1(n5462), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9108.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9109 (.I0(\i15/tx_fifo/buff[35][1] ), .I1(\i15/tx_fifo/buff[33][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9109.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9110 (.I0(\i15/tx_fifo/buff[32][1] ), .I1(\i15/tx_fifo/buff[34][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9110.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9111 (.I0(n5281), .I1(n5464), .I2(n5465), .O(n5466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9111.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9112 (.I0(\i15/tx_fifo/buff[43][1] ), .I1(\i15/tx_fifo/buff[41][1] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9112.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9113 (.I0(\i15/tx_fifo/buff[40][1] ), .I1(\i15/tx_fifo/buff[42][1] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9113.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9114 (.I0(n5277), .I1(n5467), .I2(n5468), .O(n5469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9114.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9115 (.I0(n5460), .I1(n5463), .I2(n5466), .I3(n5469), 
            .O(n5470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9115.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9116 (.I0(n5470), .I1(n5457), .I2(n5270), .I3(n5300), 
            .O(n5471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__9116.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__9117 (.I0(n5444), .I1(n5432), .I2(n5302), .I3(n5471), 
            .O(n5472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9117.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9118 (.I0(rx_en_tx_packet), .I1(\rx_d[1] ), .O(\data_to_tx_packet_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9118.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9119 (.I0(\data_to_tx_packet_reg[1] ), .I1(n5232), .O(n5473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9119.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9120 (.I0(n5472), .I1(n5419), .I2(n5361), .I3(n5473), 
            .O(\tx_fifo/n143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff70 */ ;
    defparam LUT__9120.LUTMASK = 16'hff70;
    EFX_LUT4 LUT__9121 (.I0(\i15/tx_fifo/buff[15][2] ), .I1(\i15/tx_fifo/buff[13][2] ), 
            .I2(n5252), .I3(\tx_fifo/rd_index[1] ), .O(n5474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__9121.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__9122 (.I0(\i15/tx_fifo/buff[7][2] ), .I1(\i15/tx_fifo/buff[5][2] ), 
            .I2(n5252), .I3(n5474), .O(n5475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcfa0 */ ;
    defparam LUT__9122.LUTMASK = 16'hcfa0;
    EFX_LUT4 LUT__9123 (.I0(\i15/tx_fifo/buff[3][2] ), .I1(\i15/tx_fifo/buff[1][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9123.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9124 (.I0(\i15/tx_fifo/buff[0][2] ), .I1(\i15/tx_fifo/buff[2][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9124.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9125 (.I0(\i15/tx_fifo/buff[4][2] ), .I1(\i15/tx_fifo/buff[6][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9125.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9126 (.I0(n5476), .I1(n5477), .I2(n5478), .I3(n5241), 
            .O(n5479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__9126.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__9127 (.I0(\i15/tx_fifo/buff[11][2] ), .I1(\i15/tx_fifo/buff[9][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9127.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9128 (.I0(\i15/tx_fifo/buff[8][2] ), .I1(\i15/tx_fifo/buff[10][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9128.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9129 (.I0(\i15/tx_fifo/buff[12][2] ), .I1(\i15/tx_fifo/buff[14][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9129.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9130 (.I0(n5480), .I1(n5481), .I2(n5482), .I3(n5241), 
            .O(n5483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__9130.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__9131 (.I0(n5483), .I1(n5479), .I2(n5252), .O(n5484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__9131.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__9132 (.I0(n5475), .I1(\tx_fifo/rd_index[0] ), .I2(n5241), 
            .I3(n5484), .O(n5485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9132.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9133 (.I0(\i15/tx_fifo/buff[95][2] ), .I1(\i15/tx_fifo/buff[93][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9133.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9134 (.I0(\i15/tx_fifo/buff[92][2] ), .I1(\i15/tx_fifo/buff[94][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9134.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9135 (.I0(n5486), .I1(n5487), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9135.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9136 (.I0(\i15/tx_fifo/buff[91][2] ), .I1(\i15/tx_fifo/buff[89][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9136.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9137 (.I0(\i15/tx_fifo/buff[88][2] ), .I1(\i15/tx_fifo/buff[90][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9137.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9138 (.I0(n5277), .I1(n5489), .I2(n5490), .O(n5491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9138.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9139 (.I0(\i15/tx_fifo/buff[83][2] ), .I1(\i15/tx_fifo/buff[81][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9139.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9140 (.I0(\i15/tx_fifo/buff[80][2] ), .I1(\i15/tx_fifo/buff[82][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9140.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9141 (.I0(n5281), .I1(n5492), .I2(n5493), .O(n5494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9141.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9142 (.I0(\i15/tx_fifo/buff[87][2] ), .I1(\i15/tx_fifo/buff[85][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9142.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9143 (.I0(\i15/tx_fifo/buff[84][2] ), .I1(\i15/tx_fifo/buff[86][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9143.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9144 (.I0(n5495), .I1(n5496), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9144.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9145 (.I0(n5488), .I1(n5491), .I2(n5494), .I3(n5497), 
            .O(n5498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9145.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9146 (.I0(\i15/tx_fifo/buff[79][2] ), .I1(\i15/tx_fifo/buff[77][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9146.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9147 (.I0(\i15/tx_fifo/buff[76][2] ), .I1(\i15/tx_fifo/buff[78][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9147.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9148 (.I0(n5499), .I1(n5500), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9148.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9149 (.I0(\i15/tx_fifo/buff[75][2] ), .I1(\i15/tx_fifo/buff[73][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9149.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9150 (.I0(\i15/tx_fifo/buff[72][2] ), .I1(\i15/tx_fifo/buff[74][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9150.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9151 (.I0(n5277), .I1(n5502), .I2(n5503), .O(n5504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9151.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9152 (.I0(\i15/tx_fifo/buff[67][2] ), .I1(\i15/tx_fifo/buff[65][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9152.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9153 (.I0(\i15/tx_fifo/buff[64][2] ), .I1(\i15/tx_fifo/buff[66][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9153.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9154 (.I0(n5281), .I1(n5505), .I2(n5506), .O(n5507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9154.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9155 (.I0(\i15/tx_fifo/buff[71][2] ), .I1(\i15/tx_fifo/buff[69][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9155.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9156 (.I0(\i15/tx_fifo/buff[68][2] ), .I1(\i15/tx_fifo/buff[70][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9156.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9157 (.I0(n5508), .I1(n5509), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9157.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9158 (.I0(n5501), .I1(n5504), .I2(n5507), .I3(n5510), 
            .O(n5511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9158.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9159 (.I0(n5511), .I1(n5498), .I2(n5269), .I3(n5270), 
            .O(n5512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__9159.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__9160 (.I0(\i15/tx_fifo/buff[28][2] ), .I1(\i15/tx_fifo/buff[20][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[3] ), .O(n5513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9160.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9161 (.I0(\i15/tx_fifo/buff[30][2] ), .I1(\i15/tx_fifo/buff[22][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(n5513), .O(n5514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9161.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9162 (.I0(\i15/tx_fifo/buff[31][2] ), .I1(\i15/tx_fifo/buff[29][2] ), 
            .I2(\tx_fifo/rd_index[3] ), .I3(\tx_fifo/rd_index[1] ), .O(n5515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9162.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9163 (.I0(\i15/tx_fifo/buff[21][2] ), .I1(\i15/tx_fifo/buff[23][2] ), 
            .I2(\tx_fifo/rd_index[3] ), .I3(n5515), .O(n5516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__9163.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__9164 (.I0(n5516), .I1(n5514), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9164.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9165 (.I0(\i15/tx_fifo/buff[19][2] ), .I1(\i15/tx_fifo/buff[17][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9165.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9166 (.I0(\i15/tx_fifo/buff[16][2] ), .I1(\i15/tx_fifo/buff[18][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9166.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9167 (.I0(n5518), .I1(n5519), .I2(n5281), .I3(n5270), 
            .O(n5520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9167.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9168 (.I0(\i15/tx_fifo/buff[27][2] ), .I1(\i15/tx_fifo/buff[25][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9168.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9169 (.I0(\i15/tx_fifo/buff[24][2] ), .I1(\i15/tx_fifo/buff[26][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9169.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9170 (.I0(n5521), .I1(n5522), .I2(n5277), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9170.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9171 (.I0(n5517), .I1(n5523), .I2(n5520), .I3(n5330), 
            .O(n5524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9171.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9172 (.I0(n5270), .I1(n5485), .I2(n5524), .I3(n5512), 
            .O(n5525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__9172.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__9173 (.I0(\i15/tx_fifo/buff[32][2] ), .I1(\i15/tx_fifo/buff[34][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9173.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9174 (.I0(\i15/tx_fifo/buff[35][2] ), .I1(\i15/tx_fifo/buff[33][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5526), .O(n5527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9174.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9175 (.I0(\i15/tx_fifo/buff[47][2] ), .I1(\i15/tx_fifo/buff[45][2] ), 
            .I2(\tx_fifo/rd_index[3] ), .I3(\tx_fifo/rd_index[1] ), .O(n5528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9175.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9176 (.I0(\i15/tx_fifo/buff[37][2] ), .I1(\i15/tx_fifo/buff[39][2] ), 
            .I2(\tx_fifo/rd_index[3] ), .I3(n5528), .O(n5529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__9176.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__9177 (.I0(\i15/tx_fifo/buff[44][2] ), .I1(\i15/tx_fifo/buff[46][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9177.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9178 (.I0(\i15/tx_fifo/buff[36][2] ), .I1(\i15/tx_fifo/buff[38][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9178.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9179 (.I0(n5531), .I1(n5530), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__9179.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__9180 (.I0(\i15/tx_fifo/buff[43][2] ), .I1(\i15/tx_fifo/buff[41][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9180.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9181 (.I0(\i15/tx_fifo/buff[40][2] ), .I1(\i15/tx_fifo/buff[42][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9181.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9182 (.I0(n5533), .I1(n5534), .I2(n5277), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9182.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9183 (.I0(n5529), .I1(\tx_fifo/rd_index[0] ), .I2(n5532), 
            .I3(n5535), .O(n5536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__9183.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__9184 (.I0(n5281), .I1(n5527), .I2(n5270), .I3(n5536), 
            .O(n5537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__9184.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__9185 (.I0(\i15/tx_fifo/buff[63][2] ), .I1(\i15/tx_fifo/buff[61][2] ), 
            .I2(\tx_fifo/rd_index[3] ), .I3(\tx_fifo/rd_index[1] ), .O(n5538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__9185.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__9186 (.I0(\i15/tx_fifo/buff[55][2] ), .I1(\i15/tx_fifo/buff[53][2] ), 
            .I2(\tx_fifo/rd_index[3] ), .I3(n5538), .O(n5539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__9186.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__9187 (.I0(\i15/tx_fifo/buff[52][2] ), .I1(\i15/tx_fifo/buff[54][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9187.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9188 (.I0(\i15/tx_fifo/buff[60][2] ), .I1(\i15/tx_fifo/buff[62][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9188.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9189 (.I0(n5540), .I1(n5541), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__9189.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__9190 (.I0(\i15/tx_fifo/buff[48][2] ), .I1(\i15/tx_fifo/buff[50][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9190.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9191 (.I0(\i15/tx_fifo/buff[51][2] ), .I1(\i15/tx_fifo/buff[49][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5543), .O(n5544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9191.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9192 (.I0(\i15/tx_fifo/buff[56][2] ), .I1(\i15/tx_fifo/buff[58][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9192.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9193 (.I0(\i15/tx_fifo/buff[59][2] ), .I1(\i15/tx_fifo/buff[57][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9193.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9194 (.I0(n5546), .I1(n5545), .I2(n5277), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9194.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9195 (.I0(n5281), .I1(n5544), .I2(n5547), .I3(n5270), 
            .O(n5548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__9195.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__9196 (.I0(n5539), .I1(\tx_fifo/rd_index[0] ), .I2(n5542), 
            .I3(n5548), .O(n5549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__9196.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__9197 (.I0(\i15/tx_fifo/buff[123][2] ), .I1(\i15/tx_fifo/buff[121][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9197.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9198 (.I0(\i15/tx_fifo/buff[120][2] ), .I1(\i15/tx_fifo/buff[122][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9198.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9199 (.I0(n5277), .I1(n5550), .I2(n5551), .O(n5552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9199.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9200 (.I0(\i15/tx_fifo/buff[115][2] ), .I1(\i15/tx_fifo/buff[113][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9200.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9201 (.I0(\i15/tx_fifo/buff[112][2] ), .I1(\i15/tx_fifo/buff[114][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9201.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9202 (.I0(n5281), .I1(n5553), .I2(n5554), .O(n5555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9202.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9203 (.I0(\i15/tx_fifo/buff[119][2] ), .I1(\i15/tx_fifo/buff[117][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9203.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9204 (.I0(\i15/tx_fifo/buff[116][2] ), .I1(\i15/tx_fifo/buff[118][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9204.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9205 (.I0(n5556), .I1(n5557), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9205.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9206 (.I0(\i15/tx_fifo/buff[127][2] ), .I1(\i15/tx_fifo/buff[125][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9206.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9207 (.I0(\i15/tx_fifo/buff[124][2] ), .I1(\i15/tx_fifo/buff[126][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9207.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9208 (.I0(n5559), .I1(n5560), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9208.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9209 (.I0(n5552), .I1(n5555), .I2(n5558), .I3(n5561), 
            .O(n5562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9209.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9210 (.I0(\i15/tx_fifo/buff[99][2] ), .I1(\i15/tx_fifo/buff[97][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9210.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9211 (.I0(\i15/tx_fifo/buff[96][2] ), .I1(\i15/tx_fifo/buff[98][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9211.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9212 (.I0(n5281), .I1(n5563), .I2(n5564), .O(n5565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9212.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9213 (.I0(\i15/tx_fifo/buff[104][2] ), .I1(\i15/tx_fifo/buff[106][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9213.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9214 (.I0(\i15/tx_fifo/buff[107][2] ), .I1(\i15/tx_fifo/buff[105][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9214.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9215 (.I0(n5567), .I1(n5566), .I2(n5277), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9215.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9216 (.I0(\i15/tx_fifo/buff[103][2] ), .I1(\i15/tx_fifo/buff[101][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9216.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9217 (.I0(\i15/tx_fifo/buff[100][2] ), .I1(\i15/tx_fifo/buff[102][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9217.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9218 (.I0(n5569), .I1(n5570), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9218.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9219 (.I0(\i15/tx_fifo/buff[111][2] ), .I1(\i15/tx_fifo/buff[109][2] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9219.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9220 (.I0(\i15/tx_fifo/buff[108][2] ), .I1(\i15/tx_fifo/buff[110][2] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9220.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9221 (.I0(n5572), .I1(n5573), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9221.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9222 (.I0(n5565), .I1(n5568), .I2(n5571), .I3(n5574), 
            .O(n5575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9222.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9223 (.I0(n5575), .I1(n5562), .I2(n5270), .I3(n5302), 
            .O(n5576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__9223.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__9224 (.I0(n5549), .I1(n5537), .I2(n5300), .I3(n5576), 
            .O(n5577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9224.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9225 (.I0(rx_en_tx_packet), .I1(\rx_d[2] ), .O(\data_to_tx_packet_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9225.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9226 (.I0(\data_to_tx_packet_reg[2] ), .I1(n5232), .O(n5578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9226.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9227 (.I0(n5577), .I1(n5525), .I2(n5361), .I3(n5578), 
            .O(\tx_fifo/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff70 */ ;
    defparam LUT__9227.LUTMASK = 16'hff70;
    EFX_LUT4 LUT__9228 (.I0(\i15/tx_fifo/buff[47][3] ), .I1(\i15/tx_fifo/buff[45][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9228.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9229 (.I0(\i15/tx_fifo/buff[44][3] ), .I1(\i15/tx_fifo/buff[46][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9229.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9230 (.I0(n5579), .I1(n5580), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9230.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9231 (.I0(\i15/tx_fifo/buff[40][3] ), .I1(\i15/tx_fifo/buff[42][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9231.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9232 (.I0(\i15/tx_fifo/buff[43][3] ), .I1(\i15/tx_fifo/buff[41][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9232.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9233 (.I0(n5583), .I1(n5582), .I2(n5277), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9233.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9234 (.I0(\i15/tx_fifo/buff[35][3] ), .I1(\i15/tx_fifo/buff[33][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9234.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9235 (.I0(\i15/tx_fifo/buff[32][3] ), .I1(\i15/tx_fifo/buff[34][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9235.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9236 (.I0(\i15/tx_fifo/buff[39][3] ), .I1(\i15/tx_fifo/buff[37][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9236.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9237 (.I0(\i15/tx_fifo/buff[36][3] ), .I1(\i15/tx_fifo/buff[38][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9237.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9238 (.I0(n5587), .I1(n5588), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9238.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9239 (.I0(n5585), .I1(n5586), .I2(n5281), .I3(n5589), 
            .O(n5590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9239.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9240 (.I0(n5581), .I1(n5584), .I2(n5270), .I3(n5590), 
            .O(n5591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9240.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9241 (.I0(\i15/tx_fifo/buff[48][3] ), .I1(\i15/tx_fifo/buff[50][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9241.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9242 (.I0(\i15/tx_fifo/buff[51][3] ), .I1(\i15/tx_fifo/buff[49][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5592), .O(n5593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9242.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9243 (.I0(\i15/tx_fifo/buff[55][3] ), .I1(\i15/tx_fifo/buff[53][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9243.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9244 (.I0(n5594), .I1(\tx_fifo/rd_index[3] ), .I2(n5241), 
            .O(n5595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__9244.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__9245 (.I0(\i15/tx_fifo/buff[52][3] ), .I1(\i15/tx_fifo/buff[54][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9245.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9246 (.I0(\i15/tx_fifo/buff[63][3] ), .I1(\i15/tx_fifo/buff[61][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9246.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9247 (.I0(\i15/tx_fifo/buff[60][3] ), .I1(\i15/tx_fifo/buff[62][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9247.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9248 (.I0(n5597), .I1(n5598), .I2(n5596), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__9248.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__9249 (.I0(n5599), .I1(n5595), .I2(n5593), .I3(n5281), 
            .O(n5600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0 */ ;
    defparam LUT__9249.LUTMASK = 16'hbbb0;
    EFX_LUT4 LUT__9250 (.I0(\i15/tx_fifo/buff[59][3] ), .I1(\i15/tx_fifo/buff[57][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9250.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9251 (.I0(\i15/tx_fifo/buff[56][3] ), .I1(\i15/tx_fifo/buff[58][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9251.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9252 (.I0(n5601), .I1(n5602), .I2(n5277), .I3(n5270), 
            .O(n5603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9252.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9253 (.I0(n5603), .I1(n5600), .I2(n5300), .O(n5604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__9253.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__9254 (.I0(\i15/tx_fifo/buff[111][3] ), .I1(\i15/tx_fifo/buff[109][3] ), 
            .I2(\tx_fifo/rd_index[3] ), .I3(\tx_fifo/rd_index[1] ), .O(n5605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__9254.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__9255 (.I0(\i15/tx_fifo/buff[103][3] ), .I1(\i15/tx_fifo/buff[101][3] ), 
            .I2(\tx_fifo/rd_index[3] ), .I3(n5605), .O(n5606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__9255.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__9256 (.I0(\i15/tx_fifo/buff[100][3] ), .I1(\i15/tx_fifo/buff[102][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9256.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9257 (.I0(\i15/tx_fifo/buff[108][3] ), .I1(\i15/tx_fifo/buff[110][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9257.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9258 (.I0(n5607), .I1(n5608), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__9258.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__9259 (.I0(\i15/tx_fifo/buff[104][3] ), .I1(\i15/tx_fifo/buff[106][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9259.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9260 (.I0(\i15/tx_fifo/buff[107][3] ), .I1(\i15/tx_fifo/buff[105][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5610), .O(n5611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9260.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9261 (.I0(\i15/tx_fifo/buff[96][3] ), .I1(\i15/tx_fifo/buff[98][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9261.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9262 (.I0(\i15/tx_fifo/buff[99][3] ), .I1(\i15/tx_fifo/buff[97][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9262.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9263 (.I0(n5613), .I1(n5612), .I2(n5281), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9263.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9264 (.I0(n5277), .I1(n5611), .I2(n5270), .I3(n5614), 
            .O(n5615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__9264.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__9265 (.I0(n5606), .I1(\tx_fifo/rd_index[0] ), .I2(n5609), 
            .I3(n5615), .O(n5616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__9265.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__9266 (.I0(\i15/tx_fifo/buff[112][3] ), .I1(\i15/tx_fifo/buff[114][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9266.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9267 (.I0(\i15/tx_fifo/buff[115][3] ), .I1(\i15/tx_fifo/buff[113][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5617), .O(n5618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9267.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9268 (.I0(\i15/tx_fifo/buff[119][3] ), .I1(\i15/tx_fifo/buff[117][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5619)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9268.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9269 (.I0(n5619), .I1(\tx_fifo/rd_index[3] ), .I2(n5241), 
            .O(n5620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__9269.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__9270 (.I0(\i15/tx_fifo/buff[127][3] ), .I1(\i15/tx_fifo/buff[125][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5621)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9270.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9271 (.I0(\i15/tx_fifo/buff[124][3] ), .I1(\i15/tx_fifo/buff[126][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9271.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9272 (.I0(\i15/tx_fifo/buff[116][3] ), .I1(\i15/tx_fifo/buff[118][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9272.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9273 (.I0(n5621), .I1(n5622), .I2(n5623), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__9273.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__9274 (.I0(n5624), .I1(n5620), .I2(n5618), .I3(n5281), 
            .O(n5625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0 */ ;
    defparam LUT__9274.LUTMASK = 16'hbbb0;
    EFX_LUT4 LUT__9275 (.I0(\i15/tx_fifo/buff[123][3] ), .I1(\i15/tx_fifo/buff[121][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9275.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9276 (.I0(\i15/tx_fifo/buff[120][3] ), .I1(\i15/tx_fifo/buff[122][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9276.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9277 (.I0(n5626), .I1(n5627), .I2(n5277), .I3(n5270), 
            .O(n5628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9277.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9278 (.I0(n5628), .I1(n5625), .I2(n5302), .O(n5629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__9278.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__9279 (.I0(n5616), .I1(n5629), .I2(n5591), .I3(n5604), 
            .O(n5630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__9279.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__9280 (.I0(\i15/tx_fifo/buff[67][3] ), .I1(\i15/tx_fifo/buff[65][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9280.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9281 (.I0(\i15/tx_fifo/buff[64][3] ), .I1(\i15/tx_fifo/buff[66][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9281.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9282 (.I0(n5281), .I1(n5631), .I2(n5632), .O(n5633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9282.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9283 (.I0(\i15/tx_fifo/buff[75][3] ), .I1(\i15/tx_fifo/buff[73][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9283.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9284 (.I0(\i15/tx_fifo/buff[72][3] ), .I1(\i15/tx_fifo/buff[74][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9284.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9285 (.I0(n5277), .I1(n5634), .I2(n5635), .O(n5636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9285.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9286 (.I0(\i15/tx_fifo/buff[71][3] ), .I1(\i15/tx_fifo/buff[69][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9286.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9287 (.I0(\i15/tx_fifo/buff[68][3] ), .I1(\i15/tx_fifo/buff[70][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9287.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9288 (.I0(n5637), .I1(n5638), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9288.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9289 (.I0(\i15/tx_fifo/buff[79][3] ), .I1(\i15/tx_fifo/buff[77][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5640)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9289.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9290 (.I0(\i15/tx_fifo/buff[76][3] ), .I1(\i15/tx_fifo/buff[78][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9290.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9291 (.I0(n5640), .I1(n5641), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5642)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9291.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9292 (.I0(n5633), .I1(n5636), .I2(n5639), .I3(n5642), 
            .O(n5643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9292.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9293 (.I0(\i15/tx_fifo/buff[88][3] ), .I1(\i15/tx_fifo/buff[90][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9293.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9294 (.I0(\i15/tx_fifo/buff[91][3] ), .I1(\i15/tx_fifo/buff[89][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9294.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9295 (.I0(n5645), .I1(n5644), .I2(n5277), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9295.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9296 (.I0(\i15/tx_fifo/buff[95][3] ), .I1(\i15/tx_fifo/buff[93][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9296.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9297 (.I0(\i15/tx_fifo/buff[92][3] ), .I1(\i15/tx_fifo/buff[94][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9297.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9298 (.I0(n5647), .I1(n5648), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9298.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9299 (.I0(\i15/tx_fifo/buff[87][3] ), .I1(\i15/tx_fifo/buff[85][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9299.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9300 (.I0(\i15/tx_fifo/buff[84][3] ), .I1(\i15/tx_fifo/buff[86][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9300.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9301 (.I0(n5650), .I1(n5651), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9301.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9302 (.I0(\i15/tx_fifo/buff[83][3] ), .I1(\i15/tx_fifo/buff[81][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9302.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9303 (.I0(\i15/tx_fifo/buff[80][3] ), .I1(\i15/tx_fifo/buff[82][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9303.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9304 (.I0(n5281), .I1(n5653), .I2(n5654), .O(n5655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9304.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9305 (.I0(n5646), .I1(n5649), .I2(n5652), .I3(n5655), 
            .O(n5656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9305.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9306 (.I0(n5656), .I1(n5643), .I2(n5269), .I3(n5270), 
            .O(n5657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9306.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9307 (.I0(\i15/tx_fifo/buff[19][3] ), .I1(\i15/tx_fifo/buff[17][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9307.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9308 (.I0(\i15/tx_fifo/buff[16][3] ), .I1(\i15/tx_fifo/buff[18][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9308.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9309 (.I0(n5281), .I1(n5658), .I2(n5659), .O(n5660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9309.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9310 (.I0(\i15/tx_fifo/buff[27][3] ), .I1(\i15/tx_fifo/buff[25][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9310.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9311 (.I0(\i15/tx_fifo/buff[24][3] ), .I1(\i15/tx_fifo/buff[26][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9311.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9312 (.I0(n5277), .I1(n5661), .I2(n5662), .O(n5663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9312.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9313 (.I0(\i15/tx_fifo/buff[31][3] ), .I1(\i15/tx_fifo/buff[29][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9313.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9314 (.I0(\i15/tx_fifo/buff[28][3] ), .I1(\i15/tx_fifo/buff[30][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9314.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9315 (.I0(n5664), .I1(n5665), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9315.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9316 (.I0(\i15/tx_fifo/buff[23][3] ), .I1(\i15/tx_fifo/buff[21][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9316.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9317 (.I0(\i15/tx_fifo/buff[20][3] ), .I1(\i15/tx_fifo/buff[22][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9317.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9318 (.I0(n5667), .I1(n5668), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9318.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9319 (.I0(n5660), .I1(n5663), .I2(n5666), .I3(n5669), 
            .O(n5670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9319.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9320 (.I0(\i15/tx_fifo/buff[15][3] ), .I1(\i15/tx_fifo/buff[13][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9320.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9321 (.I0(\i15/tx_fifo/buff[12][3] ), .I1(\i15/tx_fifo/buff[14][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9321.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9322 (.I0(n5671), .I1(n5672), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9322.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9323 (.I0(\i15/tx_fifo/buff[7][3] ), .I1(\i15/tx_fifo/buff[5][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9323.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9324 (.I0(\i15/tx_fifo/buff[4][3] ), .I1(\i15/tx_fifo/buff[6][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9324.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9325 (.I0(n5674), .I1(n5675), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9325.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9326 (.I0(\i15/tx_fifo/buff[3][3] ), .I1(\i15/tx_fifo/buff[1][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5677)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9326.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9327 (.I0(\i15/tx_fifo/buff[0][3] ), .I1(\i15/tx_fifo/buff[2][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9327.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9328 (.I0(n5281), .I1(n5677), .I2(n5678), .O(n5679)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9328.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9329 (.I0(\i15/tx_fifo/buff[11][3] ), .I1(\i15/tx_fifo/buff[9][3] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9329.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9330 (.I0(\i15/tx_fifo/buff[8][3] ), .I1(\i15/tx_fifo/buff[10][3] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5681)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9330.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9331 (.I0(n5277), .I1(n5680), .I2(n5681), .O(n5682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9331.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9332 (.I0(n5673), .I1(n5676), .I2(n5679), .I3(n5682), 
            .O(n5683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9332.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9333 (.I0(n5683), .I1(n5670), .I2(n5330), .I3(n5270), 
            .O(n5684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__9333.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__9334 (.I0(n5657), .I1(n5684), .O(n5685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__9334.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__9335 (.I0(rx_en_tx_packet), .I1(\rx_d[3] ), .O(\data_to_tx_packet_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9335.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9336 (.I0(\data_to_tx_packet_reg[3] ), .I1(n5232), .O(n5686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9336.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9337 (.I0(n5685), .I1(n5630), .I2(n5361), .I3(n5686), 
            .O(\tx_fifo/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff70 */ ;
    defparam LUT__9337.LUTMASK = 16'hff70;
    EFX_LUT4 LUT__9338 (.I0(\i15/tx_fifo/buff[72][4] ), .I1(\i15/tx_fifo/buff[74][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__9338.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__9339 (.I0(\i15/tx_fifo/buff[75][4] ), .I1(\i15/tx_fifo/buff[73][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5687), .O(n5688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__9339.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__9340 (.I0(\i15/tx_fifo/buff[79][4] ), .I1(\i15/tx_fifo/buff[77][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9340.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9341 (.I0(\i15/tx_fifo/buff[76][4] ), .I1(\i15/tx_fifo/buff[78][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9341.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9342 (.I0(n5689), .I1(n5690), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9342.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9343 (.I0(\i15/tx_fifo/buff[67][4] ), .I1(\i15/tx_fifo/buff[65][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9343.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9344 (.I0(\i15/tx_fifo/buff[64][4] ), .I1(\i15/tx_fifo/buff[66][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9344.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9345 (.I0(\i15/tx_fifo/buff[71][4] ), .I1(\i15/tx_fifo/buff[69][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9345.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9346 (.I0(\i15/tx_fifo/buff[68][4] ), .I1(\i15/tx_fifo/buff[70][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9346.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9347 (.I0(n5694), .I1(n5695), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9347.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9348 (.I0(n5692), .I1(n5693), .I2(n5281), .I3(n5696), 
            .O(n5697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9348.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9349 (.I0(n5688), .I1(n5277), .I2(n5691), .I3(n5697), 
            .O(n5698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__9349.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__9350 (.I0(\i15/tx_fifo/buff[83][4] ), .I1(\i15/tx_fifo/buff[81][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5699)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9350.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9351 (.I0(\i15/tx_fifo/buff[80][4] ), .I1(\i15/tx_fifo/buff[82][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5700)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9351.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9352 (.I0(\i15/tx_fifo/buff[84][4] ), .I1(\i15/tx_fifo/buff[86][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9352.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9353 (.I0(n5699), .I1(n5700), .I2(n5701), .I3(n5241), 
            .O(n5702)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__9353.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__9354 (.I0(\i15/tx_fifo/buff[87][4] ), .I1(\i15/tx_fifo/buff[85][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9354.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9355 (.I0(\i15/tx_fifo/buff[95][4] ), .I1(\i15/tx_fifo/buff[93][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9355.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9356 (.I0(\i15/tx_fifo/buff[92][4] ), .I1(\i15/tx_fifo/buff[94][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9356.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9357 (.I0(n5704), .I1(n5705), .I2(n5703), .I3(n5252), 
            .O(n5706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__9357.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__9358 (.I0(\i15/tx_fifo/buff[91][4] ), .I1(\i15/tx_fifo/buff[89][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9358.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9359 (.I0(\i15/tx_fifo/buff[88][4] ), .I1(\i15/tx_fifo/buff[90][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9359.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9360 (.I0(n5707), .I1(n5708), .I2(n5706), .I3(n5241), 
            .O(n5709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__9360.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__9361 (.I0(n5241), .I1(n5702), .I2(n5252), .I3(n5709), 
            .O(n5710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h301f */ ;
    defparam LUT__9361.LUTMASK = 16'h301f;
    EFX_LUT4 LUT__9362 (.I0(n5710), .I1(n5698), .I2(n5269), .I3(n5270), 
            .O(n5711)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__9362.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__9363 (.I0(\i15/tx_fifo/buff[43][4] ), .I1(\i15/tx_fifo/buff[41][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5712)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9363.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9364 (.I0(\i15/tx_fifo/buff[40][4] ), .I1(\i15/tx_fifo/buff[42][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9364.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9365 (.I0(\i15/tx_fifo/buff[44][4] ), .I1(\i15/tx_fifo/buff[46][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9365.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9366 (.I0(\i15/tx_fifo/buff[47][4] ), .I1(\i15/tx_fifo/buff[45][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9366.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9367 (.I0(n5715), .I1(n5714), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9367.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9368 (.I0(n5713), .I1(n5241), .I2(n5712), .I3(n5716), 
            .O(n5717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9368.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9369 (.I0(\i15/tx_fifo/buff[35][4] ), .I1(\i15/tx_fifo/buff[33][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9369.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9370 (.I0(\i15/tx_fifo/buff[32][4] ), .I1(\i15/tx_fifo/buff[34][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9370.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9371 (.I0(\i15/tx_fifo/buff[36][4] ), .I1(\i15/tx_fifo/buff[38][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9371.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9372 (.I0(\i15/tx_fifo/buff[39][4] ), .I1(\i15/tx_fifo/buff[37][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9372.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9373 (.I0(n5721), .I1(n5720), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9373.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9374 (.I0(n5719), .I1(n5241), .I2(n5718), .I3(n5722), 
            .O(n5723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9374.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9375 (.I0(n5723), .I1(n5717), .I2(n5252), .O(n5724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9375.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9376 (.I0(\i15/tx_fifo/buff[51][4] ), .I1(\i15/tx_fifo/buff[49][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9376.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9377 (.I0(\i15/tx_fifo/buff[48][4] ), .I1(\i15/tx_fifo/buff[50][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5726)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9377.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9378 (.I0(\i15/tx_fifo/buff[52][4] ), .I1(\i15/tx_fifo/buff[54][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9378.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9379 (.I0(\i15/tx_fifo/buff[55][4] ), .I1(\i15/tx_fifo/buff[53][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9379.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9380 (.I0(n5728), .I1(n5727), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9380.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9381 (.I0(n5726), .I1(n5241), .I2(n5725), .I3(n5729), 
            .O(n5730)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9381.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9382 (.I0(\i15/tx_fifo/buff[59][4] ), .I1(\i15/tx_fifo/buff[57][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9382.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9383 (.I0(\i15/tx_fifo/buff[56][4] ), .I1(\i15/tx_fifo/buff[58][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9383.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9384 (.I0(\i15/tx_fifo/buff[60][4] ), .I1(\i15/tx_fifo/buff[62][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9384.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9385 (.I0(\i15/tx_fifo/buff[63][4] ), .I1(\i15/tx_fifo/buff[61][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9385.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9386 (.I0(n5734), .I1(n5733), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9386.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9387 (.I0(n5732), .I1(n5241), .I2(n5731), .I3(n5735), 
            .O(n5736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9387.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9388 (.I0(n5736), .I1(n5730), .I2(n5252), .O(n5737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__9388.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__9389 (.I0(n5737), .I1(n5724), .I2(n5270), .I3(n5300), 
            .O(n5738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9389.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9390 (.I0(\i15/tx_fifo/buff[108][4] ), .I1(\i15/tx_fifo/buff[110][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9390.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9391 (.I0(\i15/tx_fifo/buff[111][4] ), .I1(\i15/tx_fifo/buff[109][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9391.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9392 (.I0(n5740), .I1(n5739), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9392.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9393 (.I0(\i15/tx_fifo/buff[104][4] ), .I1(\i15/tx_fifo/buff[106][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9393.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9394 (.I0(\i15/tx_fifo/buff[107][4] ), .I1(\i15/tx_fifo/buff[105][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9394.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9395 (.I0(n5743), .I1(n5742), .I2(n5241), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9395.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9396 (.I0(\i15/tx_fifo/buff[99][4] ), .I1(\i15/tx_fifo/buff[97][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9396.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9397 (.I0(\i15/tx_fifo/buff[96][4] ), .I1(\i15/tx_fifo/buff[98][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9397.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9398 (.I0(\i15/tx_fifo/buff[100][4] ), .I1(\i15/tx_fifo/buff[102][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9398.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9399 (.I0(\i15/tx_fifo/buff[103][4] ), .I1(\i15/tx_fifo/buff[101][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9399.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9400 (.I0(n5748), .I1(n5747), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9400.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9401 (.I0(n5746), .I1(n5241), .I2(n5745), .I3(n5749), 
            .O(n5750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9401.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9402 (.I0(n5744), .I1(n5741), .I2(n5750), .I3(n5252), 
            .O(n5751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__9402.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__9403 (.I0(\i15/tx_fifo/buff[23][4] ), .I1(\i15/tx_fifo/buff[21][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9403.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9404 (.I0(\i15/tx_fifo/buff[20][4] ), .I1(\i15/tx_fifo/buff[22][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9404.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9405 (.I0(n5752), .I1(n5753), .I2(n5241), .O(n5754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__9405.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__9406 (.I0(\i15/tx_fifo/buff[19][4] ), .I1(\i15/tx_fifo/buff[17][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9406.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9407 (.I0(\i15/tx_fifo/buff[16][4] ), .I1(\i15/tx_fifo/buff[18][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9407.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9408 (.I0(n5756), .I1(n5241), .I2(n5755), .I3(n5252), 
            .O(n5757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9408.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9409 (.I0(\i15/tx_fifo/buff[31][4] ), .I1(\i15/tx_fifo/buff[29][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9409.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9410 (.I0(\i15/tx_fifo/buff[28][4] ), .I1(\i15/tx_fifo/buff[30][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9410.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9411 (.I0(n5758), .I1(n5759), .I2(n5241), .O(n5760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__9411.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__9412 (.I0(\i15/tx_fifo/buff[27][4] ), .I1(\i15/tx_fifo/buff[25][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9412.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9413 (.I0(\i15/tx_fifo/buff[24][4] ), .I1(\i15/tx_fifo/buff[26][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9413.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9414 (.I0(n5762), .I1(n5241), .I2(n5761), .I3(n5252), 
            .O(n5763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9414.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9415 (.I0(n5760), .I1(n5763), .I2(n5754), .I3(n5757), 
            .O(n5764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__9415.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__9416 (.I0(\i15/tx_fifo/buff[7][4] ), .I1(\i15/tx_fifo/buff[5][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9416.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9417 (.I0(\i15/tx_fifo/buff[4][4] ), .I1(\i15/tx_fifo/buff[6][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5766)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9417.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9418 (.I0(n5765), .I1(n5766), .I2(n5241), .O(n5767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__9418.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__9419 (.I0(\i15/tx_fifo/buff[3][4] ), .I1(\i15/tx_fifo/buff[1][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9419.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9420 (.I0(\i15/tx_fifo/buff[0][4] ), .I1(\i15/tx_fifo/buff[2][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9420.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9421 (.I0(n5769), .I1(n5241), .I2(n5768), .I3(n5252), 
            .O(n5770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9421.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9422 (.I0(\i15/tx_fifo/buff[15][4] ), .I1(\i15/tx_fifo/buff[13][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9422.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9423 (.I0(\i15/tx_fifo/buff[12][4] ), .I1(\i15/tx_fifo/buff[14][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9423.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9424 (.I0(n5771), .I1(n5772), .I2(n5241), .O(n5773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__9424.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__9425 (.I0(\i15/tx_fifo/buff[11][4] ), .I1(\i15/tx_fifo/buff[9][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9425.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9426 (.I0(\i15/tx_fifo/buff[8][4] ), .I1(\i15/tx_fifo/buff[10][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9426.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9427 (.I0(n5775), .I1(n5241), .I2(n5774), .I3(n5252), 
            .O(n5776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9427.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9428 (.I0(n5773), .I1(n5776), .I2(n5767), .I3(n5770), 
            .O(n5777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__9428.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__9429 (.I0(n5777), .I1(n5764), .I2(n5330), .I3(n5270), 
            .O(n5778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__9429.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__9430 (.I0(\i15/tx_fifo/buff[127][4] ), .I1(\i15/tx_fifo/buff[125][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9430.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9431 (.I0(\i15/tx_fifo/buff[124][4] ), .I1(\i15/tx_fifo/buff[126][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9431.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9432 (.I0(n5779), .I1(n5780), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9432.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9433 (.I0(\i15/tx_fifo/buff[115][4] ), .I1(\i15/tx_fifo/buff[113][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9433.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9434 (.I0(\i15/tx_fifo/buff[112][4] ), .I1(\i15/tx_fifo/buff[114][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9434.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9435 (.I0(n5281), .I1(n5782), .I2(n5783), .O(n5784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9435.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9436 (.I0(\i15/tx_fifo/buff[119][4] ), .I1(\i15/tx_fifo/buff[117][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9436.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9437 (.I0(\i15/tx_fifo/buff[116][4] ), .I1(\i15/tx_fifo/buff[118][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9437.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9438 (.I0(n5785), .I1(n5786), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9438.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9439 (.I0(\i15/tx_fifo/buff[123][4] ), .I1(\i15/tx_fifo/buff[121][4] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9439.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9440 (.I0(\i15/tx_fifo/buff[120][4] ), .I1(\i15/tx_fifo/buff[122][4] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9440.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9441 (.I0(n5277), .I1(n5788), .I2(n5789), .O(n5790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9441.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9442 (.I0(n5781), .I1(n5784), .I2(n5787), .I3(n5790), 
            .O(n5791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9442.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9443 (.I0(n5360), .I1(n5791), .I2(n5361), .O(n5792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__9443.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__9444 (.I0(n5303), .I1(n5751), .I2(n5778), .I3(n5792), 
            .O(n5793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__9444.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__9445 (.I0(rx_en_tx_packet), .I1(\rx_d[4] ), .O(\data_to_tx_packet_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9445.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9446 (.I0(\data_to_tx_packet_reg[4] ), .I1(n5232), .O(n5794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9446.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9447 (.I0(n5738), .I1(n5711), .I2(n5793), .I3(n5794), 
            .O(\tx_fifo/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10 */ ;
    defparam LUT__9447.LUTMASK = 16'hff10;
    EFX_LUT4 LUT__9448 (.I0(\i15/tx_fifo/buff[39][5] ), .I1(\i15/tx_fifo/buff[37][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9448.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9449 (.I0(\i15/tx_fifo/buff[36][5] ), .I1(\i15/tx_fifo/buff[38][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9449.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9450 (.I0(\i15/tx_fifo/buff[32][5] ), .I1(\i15/tx_fifo/buff[34][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9450.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9451 (.I0(\i15/tx_fifo/buff[35][5] ), .I1(\i15/tx_fifo/buff[33][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5797), .O(n5798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9451.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9452 (.I0(n5796), .I1(n5795), .I2(n5798), .I3(n5241), 
            .O(n5799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__9452.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__9453 (.I0(\i15/tx_fifo/buff[43][5] ), .I1(\i15/tx_fifo/buff[41][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9453.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9454 (.I0(\i15/tx_fifo/buff[40][5] ), .I1(\i15/tx_fifo/buff[42][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9454.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9455 (.I0(\i15/tx_fifo/buff[44][5] ), .I1(\i15/tx_fifo/buff[46][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9455.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9456 (.I0(\i15/tx_fifo/buff[47][5] ), .I1(\i15/tx_fifo/buff[45][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9456.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9457 (.I0(n5803), .I1(n5802), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9457.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9458 (.I0(n5801), .I1(n5241), .I2(n5800), .I3(n5804), 
            .O(n5805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9458.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9459 (.I0(n5805), .I1(n5799), .I2(n5252), .O(n5806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__9459.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__9460 (.I0(\i15/tx_fifo/buff[59][5] ), .I1(\i15/tx_fifo/buff[57][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9460.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9461 (.I0(\i15/tx_fifo/buff[56][5] ), .I1(\i15/tx_fifo/buff[58][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9461.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9462 (.I0(\i15/tx_fifo/buff[60][5] ), .I1(\i15/tx_fifo/buff[62][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9462.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9463 (.I0(\i15/tx_fifo/buff[63][5] ), .I1(\i15/tx_fifo/buff[61][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9463.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9464 (.I0(n5810), .I1(n5809), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9464.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9465 (.I0(n5808), .I1(n5241), .I2(n5807), .I3(n5811), 
            .O(n5812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9465.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9466 (.I0(\i15/tx_fifo/buff[55][5] ), .I1(\i15/tx_fifo/buff[53][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9466.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9467 (.I0(\i15/tx_fifo/buff[52][5] ), .I1(\i15/tx_fifo/buff[54][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5814)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9467.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9468 (.I0(\i15/tx_fifo/buff[48][5] ), .I1(\i15/tx_fifo/buff[50][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9468.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9469 (.I0(\i15/tx_fifo/buff[51][5] ), .I1(\i15/tx_fifo/buff[49][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5815), .O(n5816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9469.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9470 (.I0(n5814), .I1(n5813), .I2(n5816), .I3(n5241), 
            .O(n5817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__9470.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__9471 (.I0(n5817), .I1(n5812), .I2(n5252), .O(n5818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9471.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9472 (.I0(n5818), .I1(n5806), .I2(n5270), .I3(n5300), 
            .O(n5819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__9472.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__9473 (.I0(\i15/tx_fifo/buff[95][5] ), .I1(\i15/tx_fifo/buff[93][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9473.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9474 (.I0(\i15/tx_fifo/buff[92][5] ), .I1(\i15/tx_fifo/buff[94][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9474.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9475 (.I0(\i15/tx_fifo/buff[91][5] ), .I1(\i15/tx_fifo/buff[89][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9475.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9476 (.I0(\i15/tx_fifo/buff[88][5] ), .I1(\i15/tx_fifo/buff[90][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9476.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9477 (.I0(n5822), .I1(n5823), .I2(n5821), .I3(n5241), 
            .O(n5824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__9477.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__9478 (.I0(n5820), .I1(n5241), .I2(n5252), .I3(n5824), 
            .O(n5825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0c */ ;
    defparam LUT__9478.LUTMASK = 16'h0b0c;
    EFX_LUT4 LUT__9479 (.I0(\i15/tx_fifo/buff[83][5] ), .I1(\i15/tx_fifo/buff[81][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9479.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9480 (.I0(\i15/tx_fifo/buff[80][5] ), .I1(\i15/tx_fifo/buff[82][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9480.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9481 (.I0(\i15/tx_fifo/buff[84][5] ), .I1(\i15/tx_fifo/buff[86][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9481.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9482 (.I0(n5826), .I1(n5827), .I2(n5828), .I3(n5241), 
            .O(n5829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__9482.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__9483 (.I0(\i15/tx_fifo/buff[87][5] ), .I1(\i15/tx_fifo/buff[85][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9483.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9484 (.I0(n5830), .I1(n5241), .I2(n5829), .I3(n5252), 
            .O(n5831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__9484.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__9485 (.I0(n5825), .I1(n5831), .I2(n5270), .I3(n5361), 
            .O(n5832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9485.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9486 (.I0(\i15/tx_fifo/buff[71][5] ), .I1(\i15/tx_fifo/buff[69][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9486.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9487 (.I0(\i15/tx_fifo/buff[68][5] ), .I1(\i15/tx_fifo/buff[70][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9487.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9488 (.I0(\i15/tx_fifo/buff[67][5] ), .I1(\i15/tx_fifo/buff[65][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9488.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9489 (.I0(\i15/tx_fifo/buff[64][5] ), .I1(\i15/tx_fifo/buff[66][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9489.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9490 (.I0(n5835), .I1(n5836), .I2(n5834), .I3(n5241), 
            .O(n5837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__9490.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__9491 (.I0(n5833), .I1(n5241), .I2(n5837), .I3(n5252), 
            .O(n5838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__9491.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__9492 (.I0(\i15/tx_fifo/buff[79][5] ), .I1(\i15/tx_fifo/buff[77][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9492.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9493 (.I0(\i15/tx_fifo/buff[76][5] ), .I1(\i15/tx_fifo/buff[78][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9493.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9494 (.I0(\i15/tx_fifo/buff[75][5] ), .I1(\i15/tx_fifo/buff[73][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9494.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9495 (.I0(\i15/tx_fifo/buff[72][5] ), .I1(\i15/tx_fifo/buff[74][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9495.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9496 (.I0(n5842), .I1(n5241), .I2(n5841), .I3(n5252), 
            .O(n5843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9496.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9497 (.I0(n5839), .I1(n5840), .I2(n5241), .I3(n5843), 
            .O(n5844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9497.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9498 (.I0(n5838), .I1(n5844), .I2(n5270), .I3(n5361), 
            .O(n5845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9498.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9499 (.I0(n5269), .I1(n5361), .I2(n5832), .I3(n5845), 
            .O(n5846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__9499.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__9500 (.I0(\i15/tx_fifo/buff[108][5] ), .I1(\i15/tx_fifo/buff[110][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9500.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9501 (.I0(\i15/tx_fifo/buff[111][5] ), .I1(\i15/tx_fifo/buff[109][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5847), .O(n5848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__9501.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__9502 (.I0(\i15/tx_fifo/buff[107][5] ), .I1(\i15/tx_fifo/buff[105][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9502.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9503 (.I0(\i15/tx_fifo/buff[104][5] ), .I1(\i15/tx_fifo/buff[106][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5850)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9503.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9504 (.I0(n5850), .I1(n5241), .I2(n5849), .I3(n5252), 
            .O(n5851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9504.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9505 (.I0(n5241), .I1(n5848), .I2(n5847), .I3(n5851), 
            .O(n5852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7d00 */ ;
    defparam LUT__9505.LUTMASK = 16'h7d00;
    EFX_LUT4 LUT__9506 (.I0(\i15/tx_fifo/buff[103][5] ), .I1(\i15/tx_fifo/buff[101][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9506.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9507 (.I0(\i15/tx_fifo/buff[100][5] ), .I1(\i15/tx_fifo/buff[102][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9507.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9508 (.I0(\i15/tx_fifo/buff[99][5] ), .I1(\i15/tx_fifo/buff[97][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9508.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9509 (.I0(\i15/tx_fifo/buff[96][5] ), .I1(\i15/tx_fifo/buff[98][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9509.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9510 (.I0(n5856), .I1(n5241), .I2(n5855), .I3(n5252), 
            .O(n5857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9510.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9511 (.I0(n5853), .I1(n5854), .I2(n5241), .I3(n5857), 
            .O(n5858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9511.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9512 (.I0(n5858), .I1(n5852), .I2(n5270), .I3(n5302), 
            .O(n5859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__9512.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__9513 (.I0(\i15/tx_fifo/buff[24][5] ), .I1(\i15/tx_fifo/buff[26][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9513.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9514 (.I0(\i15/tx_fifo/buff[27][5] ), .I1(\i15/tx_fifo/buff[25][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5860), .O(n5861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9514.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9515 (.I0(\i15/tx_fifo/buff[28][5] ), .I1(\i15/tx_fifo/buff[30][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9515.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9516 (.I0(\i15/tx_fifo/buff[31][5] ), .I1(\i15/tx_fifo/buff[29][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5862), .O(n5863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9516.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9517 (.I0(n5863), .I1(n5861), .I2(n5252), .I3(n5241), 
            .O(n5864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__9517.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__9518 (.I0(\i15/tx_fifo/buff[19][5] ), .I1(\i15/tx_fifo/buff[17][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9518.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9519 (.I0(\i15/tx_fifo/buff[16][5] ), .I1(\i15/tx_fifo/buff[18][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9519.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9520 (.I0(n5241), .I1(n5865), .I2(n5866), .I3(n5252), 
            .O(n5867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9520.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9521 (.I0(\i15/tx_fifo/buff[23][5] ), .I1(\i15/tx_fifo/buff[21][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9521.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9522 (.I0(\tx_fifo/rd_index[1] ), .I1(\i15/tx_fifo/buff[22][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .O(n5869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__9522.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__9523 (.I0(\tx_fifo/rd_index[2] ), .I1(\i15/tx_fifo/buff[20][5] ), 
            .O(n5870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__9523.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__9524 (.I0(n5868), .I1(n5869), .I2(n5870), .I3(n5241), 
            .O(n5871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9524.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9525 (.I0(n5871), .I1(n5867), .I2(n5864), .I3(n5331), 
            .O(n5872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__9525.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__9526 (.I0(\i15/tx_fifo/buff[127][5] ), .I1(\i15/tx_fifo/buff[125][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9526.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9527 (.I0(\i15/tx_fifo/buff[124][5] ), .I1(\i15/tx_fifo/buff[126][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9527.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9528 (.I0(\i15/tx_fifo/buff[123][5] ), .I1(\i15/tx_fifo/buff[121][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9528.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9529 (.I0(\i15/tx_fifo/buff[120][5] ), .I1(\i15/tx_fifo/buff[122][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9529.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9530 (.I0(n5875), .I1(n5876), .I2(n5241), .O(n5877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9530.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9531 (.I0(n5873), .I1(n5874), .I2(n5241), .I3(n5877), 
            .O(n5878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9531.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9532 (.I0(\i15/tx_fifo/buff[119][5] ), .I1(\i15/tx_fifo/buff[117][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9532.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9533 (.I0(\i15/tx_fifo/buff[116][5] ), .I1(\i15/tx_fifo/buff[118][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9533.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9534 (.I0(\i15/tx_fifo/buff[112][5] ), .I1(\i15/tx_fifo/buff[114][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9534.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9535 (.I0(\i15/tx_fifo/buff[115][5] ), .I1(\i15/tx_fifo/buff[113][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5881), .O(n5882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9535.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9536 (.I0(n5880), .I1(n5879), .I2(n5882), .I3(n5241), 
            .O(n5883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__9536.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__9537 (.I0(n5883), .I1(n5878), .I2(n5252), .I3(n5360), 
            .O(n5884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__9537.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__9538 (.I0(\i15/tx_fifo/buff[11][5] ), .I1(\i15/tx_fifo/buff[9][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9538.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9539 (.I0(\i15/tx_fifo/buff[8][5] ), .I1(\i15/tx_fifo/buff[10][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9539.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9540 (.I0(\i15/tx_fifo/buff[12][5] ), .I1(\i15/tx_fifo/buff[14][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9540.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9541 (.I0(\i15/tx_fifo/buff[15][5] ), .I1(\i15/tx_fifo/buff[13][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5887), .O(n5888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9541.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9542 (.I0(n5886), .I1(n5885), .I2(n5888), .I3(n5241), 
            .O(n5889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__9542.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__9543 (.I0(\i15/tx_fifo/buff[3][5] ), .I1(\i15/tx_fifo/buff[1][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9543.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9544 (.I0(\i15/tx_fifo/buff[0][5] ), .I1(\i15/tx_fifo/buff[2][5] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9544.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9545 (.I0(\i15/tx_fifo/buff[4][5] ), .I1(\i15/tx_fifo/buff[6][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9545.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9546 (.I0(\i15/tx_fifo/buff[7][5] ), .I1(\i15/tx_fifo/buff[5][5] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5892), .O(n5893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9546.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9547 (.I0(n5891), .I1(n5890), .I2(n5893), .I3(n5241), 
            .O(n5894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__9547.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__9548 (.I0(n5894), .I1(n5889), .I2(n5344), .I3(n5252), 
            .O(n5895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__9548.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__9549 (.I0(n5859), .I1(n5872), .I2(n5884), .I3(n5895), 
            .O(n5896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9549.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9550 (.I0(rx_en_tx_packet), .I1(\rx_d[5] ), .O(\data_to_tx_packet_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9550.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9551 (.I0(\data_to_tx_packet_reg[5] ), .I1(n5232), .O(n5897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9551.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9552 (.I0(n5846), .I1(n5819), .I2(n5896), .I3(n5897), 
            .O(\tx_fifo/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10 */ ;
    defparam LUT__9552.LUTMASK = 16'hff10;
    EFX_LUT4 LUT__9553 (.I0(\i15/tx_fifo/buff[75][6] ), .I1(\i15/tx_fifo/buff[73][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9553.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9554 (.I0(\i15/tx_fifo/buff[72][6] ), .I1(\i15/tx_fifo/buff[74][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9554.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9555 (.I0(\i15/tx_fifo/buff[79][6] ), .I1(\i15/tx_fifo/buff[77][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9555.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9556 (.I0(\tx_fifo/rd_index[1] ), .I1(\tx_fifo/rd_index[0] ), 
            .O(n5901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__9556.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9557 (.I0(\i15/tx_fifo/buff[78][6] ), .I1(n5901), .I2(\i15/tx_fifo/buff[76][6] ), 
            .I3(\tx_fifo/rd_index[2] ), .O(n5902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0 */ ;
    defparam LUT__9557.LUTMASK = 16'hbbb0;
    EFX_LUT4 LUT__9558 (.I0(n5900), .I1(n5902), .I2(n5241), .I3(n5270), 
            .O(n5903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__9558.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__9559 (.I0(n5899), .I1(n5898), .I2(n5241), .I3(n5903), 
            .O(n5904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__9559.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__9560 (.I0(\i15/tx_fifo/buff[88][6] ), .I1(\i15/tx_fifo/buff[90][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9560.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9561 (.I0(\i15/tx_fifo/buff[91][6] ), .I1(\i15/tx_fifo/buff[89][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9561.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9562 (.I0(n5906), .I1(n5905), .I2(n5241), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9562.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9563 (.I0(\i15/tx_fifo/buff[92][6] ), .I1(\i15/tx_fifo/buff[94][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9563.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9564 (.I0(\i15/tx_fifo/buff[95][6] ), .I1(\i15/tx_fifo/buff[93][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9564.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9565 (.I0(n5909), .I1(n5908), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9565.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9566 (.I0(n5910), .I1(n5907), .I2(n5270), .I3(n5252), 
            .O(n5911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__9566.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__9567 (.I0(\i15/tx_fifo/buff[83][6] ), .I1(\i15/tx_fifo/buff[81][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9567.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9568 (.I0(\i15/tx_fifo/buff[80][6] ), .I1(\i15/tx_fifo/buff[82][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9568.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9569 (.I0(\i15/tx_fifo/buff[84][6] ), .I1(\i15/tx_fifo/buff[86][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9569.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9570 (.I0(\i15/tx_fifo/buff[87][6] ), .I1(\i15/tx_fifo/buff[85][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5914), .O(n5915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9570.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9571 (.I0(n5913), .I1(n5912), .I2(n5915), .I3(n5241), 
            .O(n5916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__9571.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__9572 (.I0(\i15/tx_fifo/buff[71][6] ), .I1(\i15/tx_fifo/buff[69][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9572.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9573 (.I0(\i15/tx_fifo/buff[68][6] ), .I1(\i15/tx_fifo/buff[70][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9573.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9574 (.I0(\i15/tx_fifo/buff[64][6] ), .I1(\i15/tx_fifo/buff[66][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9574.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9575 (.I0(\i15/tx_fifo/buff[67][6] ), .I1(\i15/tx_fifo/buff[65][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5919), .O(n5920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9575.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9576 (.I0(n5918), .I1(n5917), .I2(n5920), .I3(n5241), 
            .O(n5921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__9576.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__9577 (.I0(n5921), .I1(n5916), .I2(n5270), .I3(n5252), 
            .O(n5922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__9577.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__9578 (.I0(n5904), .I1(n5911), .I2(n5922), .I3(n5269), 
            .O(n5923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__9578.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__9579 (.I0(\i15/tx_fifo/buff[55][6] ), .I1(\i15/tx_fifo/buff[53][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9579.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9580 (.I0(\i15/tx_fifo/buff[52][6] ), .I1(\i15/tx_fifo/buff[54][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9580.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9581 (.I0(\i15/tx_fifo/buff[51][6] ), .I1(\i15/tx_fifo/buff[49][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9581.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9582 (.I0(\i15/tx_fifo/buff[48][6] ), .I1(\i15/tx_fifo/buff[50][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9582.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9583 (.I0(n5926), .I1(n5927), .I2(n5241), .O(n5928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9583.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9584 (.I0(n5924), .I1(n5925), .I2(n5241), .I3(n5928), 
            .O(n5929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9584.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9585 (.I0(\i15/tx_fifo/buff[63][6] ), .I1(\i15/tx_fifo/buff[61][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9585.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9586 (.I0(\i15/tx_fifo/buff[60][6] ), .I1(\i15/tx_fifo/buff[62][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9586.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9587 (.I0(\i15/tx_fifo/buff[56][6] ), .I1(\i15/tx_fifo/buff[58][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9587.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9588 (.I0(\i15/tx_fifo/buff[59][6] ), .I1(\i15/tx_fifo/buff[57][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5932), .O(n5933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9588.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9589 (.I0(n5931), .I1(n5930), .I2(n5933), .I3(n5241), 
            .O(n5934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__9589.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__9590 (.I0(n5934), .I1(n5929), .I2(n5252), .I3(n5270), 
            .O(n5935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__9590.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__9591 (.I0(\i15/tx_fifo/buff[32][6] ), .I1(\i15/tx_fifo/buff[34][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__9591.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__9592 (.I0(\i15/tx_fifo/buff[35][6] ), .I1(\i15/tx_fifo/buff[33][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5936), .O(n5937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__9592.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__9593 (.I0(\i15/tx_fifo/buff[38][6] ), .I1(n5901), .I2(\i15/tx_fifo/buff[36][6] ), 
            .I3(\tx_fifo/rd_index[2] ), .O(n5938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0 */ ;
    defparam LUT__9593.LUTMASK = 16'hbbb0;
    EFX_LUT4 LUT__9594 (.I0(\i15/tx_fifo/buff[39][6] ), .I1(\i15/tx_fifo/buff[37][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9594.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9595 (.I0(n5939), .I1(n5938), .I2(n5937), .I3(n5241), 
            .O(n5940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__9595.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__9596 (.I0(\i15/tx_fifo/buff[43][6] ), .I1(\i15/tx_fifo/buff[41][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9596.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9597 (.I0(\i15/tx_fifo/buff[40][6] ), .I1(\i15/tx_fifo/buff[42][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9597.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9598 (.I0(\i15/tx_fifo/buff[44][6] ), .I1(\i15/tx_fifo/buff[46][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9598.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9599 (.I0(\i15/tx_fifo/buff[47][6] ), .I1(\i15/tx_fifo/buff[45][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5943), .O(n5944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9599.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9600 (.I0(n5942), .I1(n5941), .I2(n5944), .I3(n5241), 
            .O(n5945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__9600.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__9601 (.I0(n5945), .I1(n5940), .I2(n5270), .I3(n5252), 
            .O(n5946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__9601.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__9602 (.I0(n5946), .I1(n5935), .I2(n5300), .I3(n5361), 
            .O(n5947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__9602.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__9603 (.I0(\i15/tx_fifo/buff[28][6] ), .I1(\i15/tx_fifo/buff[30][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9603.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9604 (.I0(\i15/tx_fifo/buff[31][6] ), .I1(\i15/tx_fifo/buff[29][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9604.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9605 (.I0(n5949), .I1(n5948), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n5950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9605.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9606 (.I0(\i15/tx_fifo/buff[24][6] ), .I1(\i15/tx_fifo/buff[26][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9606.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9607 (.I0(\i15/tx_fifo/buff[27][6] ), .I1(\i15/tx_fifo/buff[25][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n5952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9607.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9608 (.I0(n5952), .I1(n5951), .I2(n5241), .I3(\tx_fifo/rd_index[0] ), 
            .O(n5953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9608.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9609 (.I0(\i15/tx_fifo/buff[15][6] ), .I1(\i15/tx_fifo/buff[13][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9609.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9610 (.I0(\i15/tx_fifo/buff[12][6] ), .I1(\i15/tx_fifo/buff[14][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9610.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9611 (.I0(n5954), .I1(n5955), .I2(n5241), .O(n5956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__9611.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__9612 (.I0(\i15/tx_fifo/buff[11][6] ), .I1(\i15/tx_fifo/buff[9][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9612.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9613 (.I0(\i15/tx_fifo/buff[8][6] ), .I1(\i15/tx_fifo/buff[10][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9613.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9614 (.I0(n5957), .I1(n5958), .I2(n5241), .O(n5959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9614.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9615 (.I0(n5959), .I1(n5270), .I2(n5956), .I3(n5252), 
            .O(n5960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9615.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9616 (.I0(n5950), .I1(n5953), .I2(n5270), .I3(n5960), 
            .O(n5961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9616.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9617 (.I0(\i15/tx_fifo/buff[19][6] ), .I1(\i15/tx_fifo/buff[17][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9617.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9618 (.I0(\i15/tx_fifo/buff[16][6] ), .I1(\i15/tx_fifo/buff[18][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9618.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9619 (.I0(\i15/tx_fifo/buff[20][6] ), .I1(\i15/tx_fifo/buff[22][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9619.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9620 (.I0(n5962), .I1(n5963), .I2(n5964), .I3(n5241), 
            .O(n5965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__9620.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__9621 (.I0(\i15/tx_fifo/buff[23][6] ), .I1(\i15/tx_fifo/buff[21][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9621.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9622 (.I0(n5966), .I1(n5241), .I2(n5965), .I3(n5270), 
            .O(n5967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__9622.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__9623 (.I0(\i15/tx_fifo/buff[3][6] ), .I1(\i15/tx_fifo/buff[1][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9623.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9624 (.I0(\i15/tx_fifo/buff[0][6] ), .I1(\i15/tx_fifo/buff[2][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9624.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9625 (.I0(\i15/tx_fifo/buff[4][6] ), .I1(\i15/tx_fifo/buff[6][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9625.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9626 (.I0(n5968), .I1(n5969), .I2(n5970), .I3(n5241), 
            .O(n5971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__9626.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__9627 (.I0(\i15/tx_fifo/buff[7][6] ), .I1(\i15/tx_fifo/buff[5][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9627.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9628 (.I0(n5972), .I1(n5241), .I2(n5344), .I3(n5971), 
            .O(n5973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0c */ ;
    defparam LUT__9628.LUTMASK = 16'h0b0c;
    EFX_LUT4 LUT__9629 (.I0(n5967), .I1(n5252), .I2(n5330), .I3(n5973), 
            .O(n5974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__9629.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__9630 (.I0(\i15/tx_fifo/buff[119][6] ), .I1(\i15/tx_fifo/buff[117][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9630.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9631 (.I0(\i15/tx_fifo/buff[116][6] ), .I1(\i15/tx_fifo/buff[118][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9631.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9632 (.I0(\i15/tx_fifo/buff[115][6] ), .I1(\i15/tx_fifo/buff[113][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9632.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9633 (.I0(\i15/tx_fifo/buff[112][6] ), .I1(\i15/tx_fifo/buff[114][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9633.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9634 (.I0(n5977), .I1(n5978), .I2(n5241), .O(n5979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9634.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9635 (.I0(n5975), .I1(n5976), .I2(n5241), .I3(n5979), 
            .O(n5980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9635.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9636 (.I0(\i15/tx_fifo/buff[127][6] ), .I1(\i15/tx_fifo/buff[125][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5981)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9636.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9637 (.I0(\i15/tx_fifo/buff[124][6] ), .I1(\i15/tx_fifo/buff[126][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9637.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9638 (.I0(\i15/tx_fifo/buff[120][6] ), .I1(\i15/tx_fifo/buff[122][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9638.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9639 (.I0(\i15/tx_fifo/buff[123][6] ), .I1(\i15/tx_fifo/buff[121][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5983), .O(n5984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9639.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9640 (.I0(n5982), .I1(n5981), .I2(n5984), .I3(n5241), 
            .O(n5985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__9640.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__9641 (.I0(n5985), .I1(n5980), .I2(n5252), .I3(n5360), 
            .O(n5986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__9641.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__9642 (.I0(\i15/tx_fifo/buff[104][6] ), .I1(\i15/tx_fifo/buff[106][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9642.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9643 (.I0(\i15/tx_fifo/buff[107][6] ), .I1(\i15/tx_fifo/buff[105][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n5987), .O(n5988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9643.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9644 (.I0(\i15/tx_fifo/buff[103][6] ), .I1(\i15/tx_fifo/buff[101][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9644.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9645 (.I0(\i15/tx_fifo/buff[100][6] ), .I1(\i15/tx_fifo/buff[102][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9645.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9646 (.I0(n5989), .I1(n5990), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n5991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9646.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9647 (.I0(\i15/tx_fifo/buff[99][6] ), .I1(\i15/tx_fifo/buff[97][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9647.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9648 (.I0(\i15/tx_fifo/buff[96][6] ), .I1(\i15/tx_fifo/buff[98][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9648.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9649 (.I0(n5281), .I1(n5992), .I2(n5993), .O(n5994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9649.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9650 (.I0(\i15/tx_fifo/buff[111][6] ), .I1(\i15/tx_fifo/buff[109][6] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n5995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9650.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9651 (.I0(\i15/tx_fifo/buff[108][6] ), .I1(\i15/tx_fifo/buff[110][6] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n5996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9651.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9652 (.I0(n5995), .I1(n5996), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n5997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9652.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9653 (.I0(n5270), .I1(n5991), .I2(n5994), .I3(n5997), 
            .O(n5998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__9653.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__9654 (.I0(n5277), .I1(n5988), .I2(n5998), .I3(n5302), 
            .O(n5999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__9654.LUTMASK = 16'he000;
    EFX_LUT4 LUT__9655 (.I0(n5974), .I1(n5961), .I2(n5986), .I3(n5999), 
            .O(n6000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__9655.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__9656 (.I0(rx_en_tx_packet), .I1(\rx_d[6] ), .O(\data_to_tx_packet_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9656.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9657 (.I0(\data_to_tx_packet_reg[6] ), .I1(n5232), .O(n6001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9657.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9658 (.I0(n5923), .I1(n6000), .I2(n5947), .I3(n6001), 
            .O(\tx_fifo/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40 */ ;
    defparam LUT__9658.LUTMASK = 16'hff40;
    EFX_LUT4 LUT__9659 (.I0(\i15/tx_fifo/buff[47][7] ), .I1(\i15/tx_fifo/buff[45][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9659.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9660 (.I0(\i15/tx_fifo/buff[44][7] ), .I1(\i15/tx_fifo/buff[46][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9660.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9661 (.I0(n6002), .I1(n6003), .I2(n5241), .I3(\tx_fifo/rd_index[3] ), 
            .O(n6004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9661.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9662 (.I0(\i15/tx_fifo/buff[39][7] ), .I1(\i15/tx_fifo/buff[37][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9662.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9663 (.I0(\i15/tx_fifo/buff[36][7] ), .I1(\i15/tx_fifo/buff[38][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9663.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9664 (.I0(n6005), .I1(n6006), .I2(\tx_fifo/rd_index[3] ), 
            .I3(n5241), .O(n6007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9664.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9665 (.I0(\i15/tx_fifo/buff[43][7] ), .I1(\i15/tx_fifo/buff[41][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9665.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9666 (.I0(\i15/tx_fifo/buff[40][7] ), .I1(\i15/tx_fifo/buff[42][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9666.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9667 (.I0(\i15/tx_fifo/buff[35][7] ), .I1(\i15/tx_fifo/buff[33][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9667.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9668 (.I0(\i15/tx_fifo/buff[32][7] ), .I1(\i15/tx_fifo/buff[34][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9668.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9669 (.I0(n5281), .I1(n6010), .I2(n6011), .O(n6012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9669.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9670 (.I0(n6008), .I1(n6009), .I2(n5277), .I3(n6012), 
            .O(n6013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9670.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9671 (.I0(n6007), .I1(n6004), .I2(n6013), .I3(n5270), 
            .O(n6014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9671.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9672 (.I0(\i15/tx_fifo/buff[51][7] ), .I1(\i15/tx_fifo/buff[49][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9672.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9673 (.I0(\i15/tx_fifo/buff[48][7] ), .I1(\i15/tx_fifo/buff[50][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9673.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9674 (.I0(\i15/tx_fifo/buff[52][7] ), .I1(\i15/tx_fifo/buff[54][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n6017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9674.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9675 (.I0(\i15/tx_fifo/buff[55][7] ), .I1(\i15/tx_fifo/buff[53][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n6018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9675.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9676 (.I0(n6018), .I1(n6017), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n6019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9676.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9677 (.I0(n6016), .I1(n5241), .I2(n6015), .I3(n6019), 
            .O(n6020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9677.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9678 (.I0(\i15/tx_fifo/buff[59][7] ), .I1(\i15/tx_fifo/buff[57][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9678.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9679 (.I0(\i15/tx_fifo/buff[56][7] ), .I1(\i15/tx_fifo/buff[58][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9679.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9680 (.I0(\i15/tx_fifo/buff[60][7] ), .I1(\i15/tx_fifo/buff[62][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n6023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9680.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9681 (.I0(\i15/tx_fifo/buff[63][7] ), .I1(\i15/tx_fifo/buff[61][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n6024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9681.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9682 (.I0(n6024), .I1(n6023), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n6025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9682.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9683 (.I0(n6022), .I1(n5241), .I2(n6021), .I3(n6025), 
            .O(n6026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9683.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9684 (.I0(n6026), .I1(n6020), .I2(n5252), .I3(n5270), 
            .O(n6027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__9684.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__9685 (.I0(n6014), .I1(n6027), .I2(n5300), .O(n6028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__9685.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__9686 (.I0(\i15/tx_fifo/buff[84][7] ), .I1(\i15/tx_fifo/buff[86][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n6029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9686.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9687 (.I0(\i15/tx_fifo/buff[87][7] ), .I1(\i15/tx_fifo/buff[85][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n6030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9687.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9688 (.I0(n6030), .I1(n6029), .I2(\tx_fifo/rd_index[0] ), 
            .I3(n5241), .O(n6031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__9688.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__9689 (.I0(\i15/tx_fifo/buff[80][7] ), .I1(\i15/tx_fifo/buff[82][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n6032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9689.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9690 (.I0(\i15/tx_fifo/buff[83][7] ), .I1(\i15/tx_fifo/buff[81][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n6033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9690.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9691 (.I0(n6033), .I1(n6032), .I2(n5241), .I3(\tx_fifo/rd_index[0] ), 
            .O(n6034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9691.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9692 (.I0(n6034), .I1(n6031), .I2(n5252), .I3(n5270), 
            .O(n6035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9692.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9693 (.I0(\i15/tx_fifo/buff[95][7] ), .I1(\i15/tx_fifo/buff[93][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9693.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9694 (.I0(\i15/tx_fifo/buff[92][7] ), .I1(\i15/tx_fifo/buff[94][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9694.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9695 (.I0(\i15/tx_fifo/buff[91][7] ), .I1(\i15/tx_fifo/buff[89][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9695.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9696 (.I0(\i15/tx_fifo/buff[88][7] ), .I1(\i15/tx_fifo/buff[90][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9696.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9697 (.I0(n6039), .I1(n5241), .I2(n6038), .I3(n5252), 
            .O(n6040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9697.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9698 (.I0(n6036), .I1(n6037), .I2(n5241), .I3(n6040), 
            .O(n6041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9698.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9699 (.I0(\i15/tx_fifo/buff[68][7] ), .I1(\i15/tx_fifo/buff[70][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9699.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9700 (.I0(\i15/tx_fifo/buff[67][7] ), .I1(\i15/tx_fifo/buff[65][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9700.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9701 (.I0(\i15/tx_fifo/buff[64][7] ), .I1(\i15/tx_fifo/buff[66][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9701.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9702 (.I0(n6043), .I1(n6044), .I2(n6042), .I3(n5241), 
            .O(n6045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__9702.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__9703 (.I0(n6045), .I1(n5252), .I2(n5270), .O(n6046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__9703.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__9704 (.I0(\i15/tx_fifo/buff[75][7] ), .I1(\i15/tx_fifo/buff[73][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9704.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9705 (.I0(\i15/tx_fifo/buff[72][7] ), .I1(\i15/tx_fifo/buff[74][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9705.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9706 (.I0(\i15/tx_fifo/buff[79][7] ), .I1(\i15/tx_fifo/buff[77][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9706.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9707 (.I0(\i15/tx_fifo/buff[76][7] ), .I1(\i15/tx_fifo/buff[78][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9707.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9708 (.I0(\i15/tx_fifo/buff[71][7] ), .I1(\i15/tx_fifo/buff[69][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9708.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9709 (.I0(n6049), .I1(n6050), .I2(n6051), .I3(n5252), 
            .O(n6052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__9709.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__9710 (.I0(n6047), .I1(n6048), .I2(n6052), .I3(n5241), 
            .O(n6053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__9710.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__9711 (.I0(n5241), .I1(n5252), .I2(n6053), .I3(n6046), 
            .O(n6054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc700 */ ;
    defparam LUT__9711.LUTMASK = 16'hc700;
    EFX_LUT4 LUT__9712 (.I0(n6041), .I1(n6035), .I2(n6054), .I3(n5269), 
            .O(n6055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__9712.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__9713 (.I0(\i15/tx_fifo/buff[31][7] ), .I1(\i15/tx_fifo/buff[29][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9713.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9714 (.I0(\i15/tx_fifo/buff[28][7] ), .I1(\i15/tx_fifo/buff[30][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9714.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9715 (.I0(\i15/tx_fifo/buff[20][7] ), .I1(\i15/tx_fifo/buff[22][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9715.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9716 (.I0(\i15/tx_fifo/buff[23][7] ), .I1(\i15/tx_fifo/buff[21][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n6058), .O(n6059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9716.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9717 (.I0(n6056), .I1(n6057), .I2(n6059), .I3(\tx_fifo/rd_index[3] ), 
            .O(n6060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__9717.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__9718 (.I0(\i15/tx_fifo/buff[19][7] ), .I1(\i15/tx_fifo/buff[17][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9718.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9719 (.I0(\i15/tx_fifo/buff[16][7] ), .I1(\i15/tx_fifo/buff[18][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9719.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9720 (.I0(\i15/tx_fifo/buff[24][7] ), .I1(\i15/tx_fifo/buff[26][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n6063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9720.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9721 (.I0(\i15/tx_fifo/buff[27][7] ), .I1(\i15/tx_fifo/buff[25][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n6064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9721.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9722 (.I0(n6064), .I1(n6063), .I2(n5277), .I3(\tx_fifo/rd_index[0] ), 
            .O(n6065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9722.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9723 (.I0(n6061), .I1(n6062), .I2(n5281), .I3(n6065), 
            .O(n6066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9723.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9724 (.I0(n5241), .I1(n6060), .I2(n6066), .I3(n5331), 
            .O(n6067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__9724.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__9725 (.I0(\i15/tx_fifo/buff[7][7] ), .I1(\i15/tx_fifo/buff[5][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9725.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9726 (.I0(\i15/tx_fifo/buff[4][7] ), .I1(\i15/tx_fifo/buff[6][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9726.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9727 (.I0(\i15/tx_fifo/buff[3][7] ), .I1(\i15/tx_fifo/buff[1][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9727.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9728 (.I0(\i15/tx_fifo/buff[0][7] ), .I1(\i15/tx_fifo/buff[2][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9728.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9729 (.I0(n6070), .I1(n6071), .I2(n5241), .O(n6072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9729.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9730 (.I0(n6068), .I1(n6069), .I2(n5241), .I3(n6072), 
            .O(n6073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9730.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9731 (.I0(\i15/tx_fifo/buff[15][7] ), .I1(\i15/tx_fifo/buff[13][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9731.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9732 (.I0(\i15/tx_fifo/buff[12][7] ), .I1(\i15/tx_fifo/buff[14][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9732.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9733 (.I0(\i15/tx_fifo/buff[8][7] ), .I1(\i15/tx_fifo/buff[10][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9733.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9734 (.I0(\i15/tx_fifo/buff[11][7] ), .I1(\i15/tx_fifo/buff[9][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(n6076), .O(n6077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9734.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9735 (.I0(n6075), .I1(n6074), .I2(n6077), .I3(n5241), 
            .O(n6078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__9735.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__9736 (.I0(n6078), .I1(n6073), .I2(n5344), .I3(n5252), 
            .O(n6079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__9736.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__9737 (.I0(\i15/tx_fifo/buff[123][7] ), .I1(\i15/tx_fifo/buff[121][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9737.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9738 (.I0(\i15/tx_fifo/buff[120][7] ), .I1(\i15/tx_fifo/buff[122][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9738.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9739 (.I0(n6080), .I1(n6081), .I2(n5241), .O(n6082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9739.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9740 (.I0(\i15/tx_fifo/buff[127][7] ), .I1(\i15/tx_fifo/buff[125][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9740.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9741 (.I0(\i15/tx_fifo/buff[124][7] ), .I1(\i15/tx_fifo/buff[126][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9741.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9742 (.I0(n6083), .I1(n6084), .I2(n5241), .I3(n5252), 
            .O(n6085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9742.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9743 (.I0(\i15/tx_fifo/buff[119][7] ), .I1(\i15/tx_fifo/buff[117][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9743.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9744 (.I0(\i15/tx_fifo/buff[116][7] ), .I1(\i15/tx_fifo/buff[118][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9744.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9745 (.I0(n6086), .I1(n6087), .I2(n5241), .O(n6088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__9745.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__9746 (.I0(\i15/tx_fifo/buff[115][7] ), .I1(\i15/tx_fifo/buff[113][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9746.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9747 (.I0(\i15/tx_fifo/buff[112][7] ), .I1(\i15/tx_fifo/buff[114][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9747.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9748 (.I0(n6090), .I1(n5241), .I2(n6089), .I3(n5252), 
            .O(n6091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9748.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9749 (.I0(n6088), .I1(n6091), .I2(n6082), .I3(n6085), 
            .O(n6092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__9749.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__9750 (.I0(\i15/tx_fifo/buff[104][7] ), .I1(\i15/tx_fifo/buff[106][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n6093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9750.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9751 (.I0(\i15/tx_fifo/buff[107][7] ), .I1(\i15/tx_fifo/buff[105][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .O(n6094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__9751.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__9752 (.I0(n6094), .I1(n6093), .I2(n5241), .I3(\tx_fifo/rd_index[0] ), 
            .O(n6095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__9752.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__9753 (.I0(\i15/tx_fifo/buff[111][7] ), .I1(\i15/tx_fifo/buff[109][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9753.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9754 (.I0(\i15/tx_fifo/buff[108][7] ), .I1(\i15/tx_fifo/buff[110][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9754.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9755 (.I0(n6096), .I1(n6097), .I2(n5241), .I3(n5252), 
            .O(n6098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9755.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9756 (.I0(\i15/tx_fifo/buff[103][7] ), .I1(\i15/tx_fifo/buff[101][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9756.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9757 (.I0(\i15/tx_fifo/buff[100][7] ), .I1(\i15/tx_fifo/buff[102][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9757.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9758 (.I0(n6099), .I1(n6100), .I2(n5241), .O(n6101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__9758.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__9759 (.I0(\i15/tx_fifo/buff[99][7] ), .I1(\i15/tx_fifo/buff[97][7] ), 
            .I2(\tx_fifo/rd_index[0] ), .I3(\tx_fifo/rd_index[1] ), .O(n6102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9759.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9760 (.I0(\i15/tx_fifo/buff[96][7] ), .I1(\i15/tx_fifo/buff[98][7] ), 
            .I2(\tx_fifo/rd_index[1] ), .I3(\tx_fifo/rd_index[0] ), .O(n6103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9760.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9761 (.I0(n6103), .I1(n5241), .I2(n6102), .I3(n5252), 
            .O(n6104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9761.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9762 (.I0(n6101), .I1(n6104), .I2(n6095), .I3(n6098), 
            .O(n6105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__9762.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__9763 (.I0(n6105), .I1(n6092), .I2(n5270), .I3(n5302), 
            .O(n6106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__9763.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__9764 (.I0(n6067), .I1(n6079), .I2(n6106), .I3(n5361), 
            .O(n6107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9764.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9765 (.I0(rx_en_tx_packet), .I1(\rx_d[7] ), .O(\data_to_tx_packet_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9765.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9766 (.I0(\data_to_tx_packet_reg[7] ), .I1(n5232), .O(n6108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9766.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9767 (.I0(n6055), .I1(n6028), .I2(n6107), .I3(n6108), 
            .O(\tx_fifo/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10 */ ;
    defparam LUT__9767.LUTMASK = 16'hff10;
    EFX_LUT4 LUT__9768 (.I0(n4248), .I1(n4318), .O(rx_en_rx_packet_len)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9768.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9769 (.I0(rx_en_rx_packet_len), .I1(\rx_fifo/wr_index[0] ), 
            .O(\rx_fifo/n153 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__9769.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__9770 (.I0(\rx_fifo/sync_wr[1] ), .I1(\rx_fifo/sync_wr[0] ), 
            .O(n6109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__9770.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9771 (.I0(n4318), .I1(n4239), .I2(n4247), .I3(n6109), 
            .O(ceg_net322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__9771.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__9772 (.I0(rx_en_rx_packet_len), .I1(\rx_fifo/rd_index[0] ), 
            .O(\rx_fifo/n162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__9772.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__9773 (.I0(\rx_fifo/wr_index[2] ), .I1(\rx_fifo/rd_index[2] ), 
            .I2(\rx_fifo/wr_index[3] ), .I3(\rx_fifo/rd_index[3] ), .O(n6110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__9773.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__9774 (.I0(\rx_fifo/wr_index[6] ), .I1(\rx_fifo/rd_index[6] ), 
            .I2(\rx_fifo/wr_index[7] ), .I3(\rx_fifo/rd_index[7] ), .O(n6111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__9774.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__9775 (.I0(\rx_fifo/wr_index[0] ), .I1(\rx_fifo/rd_index[0] ), 
            .I2(\rx_fifo/wr_index[1] ), .I3(\rx_fifo/rd_index[1] ), .O(n6112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__9775.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__9776 (.I0(\rx_fifo/wr_index[4] ), .I1(\rx_fifo/rd_index[4] ), 
            .I2(\rx_fifo/wr_index[5] ), .I3(\rx_fifo/rd_index[5] ), .O(n6113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__9776.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__9777 (.I0(n6110), .I1(n6111), .I2(n6112), .I3(n6113), 
            .O(n6114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__9777.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__9778 (.I0(n6109), .I1(\rx_fifo/sync_rd[0] ), .I2(\rx_fifo/sync_rd[1] ), 
            .O(n6115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__9778.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__9779 (.I0(n6115), .I1(n6114), .I2(rx_en_rx_packet_len), 
            .O(ceg_net340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__9779.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__9780 (.I0(rx_en_rx_packet_len), .I1(\rx_d[0] ), .O(\data_to_rx_packet_len_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9780.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9781 (.I0(n4248), .I1(n4343), .O(rx_en_rx_packet)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9781.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9782 (.I0(\rx_fifo/rd_index[0] ), .I1(\rx_fifo/rd_index[1] ), 
            .I2(\rx_fifo/rd_index[2] ), .I3(\rx_fifo/rd_index[3] ), .O(n6116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__9782.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__9783 (.I0(n6116), .I1(\rx_fifo/rd_index[4] ), .I2(\rx_fifo/rd_index[5] ), 
            .O(n6117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__9783.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__9784 (.I0(n6116), .I1(\rx_fifo/rd_index[4] ), .I2(\rx_fifo/rd_index[5] ), 
            .I3(\rx_fifo/rd_index[6] ), .O(n6118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__9784.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__9785 (.I0(n6114), .I1(n6117), .I2(n6118), .I3(ceg_net322), 
            .O(n6119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9785.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9786 (.I0(\i16/rx_fifo/buff[24][0] ), .I1(\i16/rx_fifo/buff[26][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9786.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9787 (.I0(\i16/rx_fifo/buff[25][0] ), .I1(\i16/rx_fifo/buff[27][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6120), .O(n6121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__9787.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__9788 (.I0(\rx_fifo/rd_index[0] ), .I1(\rx_fifo/rd_index[1] ), 
            .I2(\rx_fifo/rd_index[2] ), .O(n6122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__9788.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__9789 (.I0(\rx_fifo/rd_index[0] ), .I1(\rx_fifo/rd_index[1] ), 
            .I2(\rx_fifo/rd_index[2] ), .I3(\rx_fifo/rd_index[3] ), .O(n6123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__9789.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__9790 (.I0(\i16/rx_fifo/buff[28][0] ), .I1(\i16/rx_fifo/buff[30][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9790.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9791 (.I0(\i16/rx_fifo/buff[31][0] ), .I1(\i16/rx_fifo/buff[29][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6124), .O(n6125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9791.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9792 (.I0(n6125), .I1(n6121), .I2(n6122), .I3(n6123), 
            .O(n6126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha300 */ ;
    defparam LUT__9792.LUTMASK = 16'ha300;
    EFX_LUT4 LUT__9793 (.I0(n6116), .I1(\rx_fifo/rd_index[4] ), .O(n6127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__9793.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__9794 (.I0(\i16/rx_fifo/buff[3][0] ), .I1(\i16/rx_fifo/buff[1][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9794.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9795 (.I0(\i16/rx_fifo/buff[0][0] ), .I1(\i16/rx_fifo/buff[2][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9795.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9796 (.I0(\i16/rx_fifo/buff[4][0] ), .I1(\i16/rx_fifo/buff[6][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .O(n6130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9796.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9797 (.I0(\i16/rx_fifo/buff[7][0] ), .I1(\i16/rx_fifo/buff[5][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .O(n6131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9797.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9798 (.I0(n6131), .I1(n6130), .I2(\rx_fifo/rd_index[0] ), 
            .I3(n6122), .O(n6132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__9798.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__9799 (.I0(n6129), .I1(n6122), .I2(n6128), .I3(n6132), 
            .O(n6133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9799.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9800 (.I0(\i16/rx_fifo/buff[11][0] ), .I1(\i16/rx_fifo/buff[9][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9800.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9801 (.I0(\i16/rx_fifo/buff[8][0] ), .I1(\i16/rx_fifo/buff[10][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9801.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9802 (.I0(\i16/rx_fifo/buff[12][0] ), .I1(\i16/rx_fifo/buff[14][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .O(n6136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9802.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9803 (.I0(\i16/rx_fifo/buff[15][0] ), .I1(\i16/rx_fifo/buff[13][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .O(n6137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9803.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9804 (.I0(n6137), .I1(n6136), .I2(\rx_fifo/rd_index[0] ), 
            .I3(n6122), .O(n6138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__9804.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__9805 (.I0(n6135), .I1(n6122), .I2(n6134), .I3(n6138), 
            .O(n6139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9805.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9806 (.I0(n6139), .I1(n6133), .I2(n6123), .O(n6140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__9806.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__9807 (.I0(\i16/rx_fifo/buff[16][0] ), .I1(\i16/rx_fifo/buff[18][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__9807.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__9808 (.I0(\i16/rx_fifo/buff[19][0] ), .I1(\i16/rx_fifo/buff[17][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6141), .O(n6142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__9808.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__9809 (.I0(\i16/rx_fifo/buff[23][0] ), .I1(\i16/rx_fifo/buff[21][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9809.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9810 (.I0(\rx_fifo/rd_index[1] ), .I1(\i16/rx_fifo/buff[22][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .O(n6144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__9810.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__9811 (.I0(\rx_fifo/rd_index[2] ), .I1(\i16/rx_fifo/buff[20][0] ), 
            .I2(n6143), .I3(n6144), .O(n6145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__9811.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__9812 (.I0(n6145), .I1(n6142), .I2(n6123), .I3(n6122), 
            .O(n6146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9812.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9813 (.I0(n6126), .I1(n6146), .I2(n6140), .I3(n6127), 
            .O(n6147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__9813.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__9814 (.I0(\i16/rx_fifo/buff[71][0] ), .I1(\i16/rx_fifo/buff[69][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9814.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9815 (.I0(\i16/rx_fifo/buff[68][0] ), .I1(\i16/rx_fifo/buff[70][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9815.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9816 (.I0(\i16/rx_fifo/buff[64][0] ), .I1(\i16/rx_fifo/buff[66][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9816.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9817 (.I0(\i16/rx_fifo/buff[67][0] ), .I1(\i16/rx_fifo/buff[65][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6150), .O(n6151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9817.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9818 (.I0(n6149), .I1(n6148), .I2(n6151), .I3(n6122), 
            .O(n6152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__9818.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__9819 (.I0(\i16/rx_fifo/buff[79][0] ), .I1(\i16/rx_fifo/buff[77][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9819.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9820 (.I0(\i16/rx_fifo/buff[76][0] ), .I1(\i16/rx_fifo/buff[78][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9820.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9821 (.I0(\i16/rx_fifo/buff[75][0] ), .I1(\i16/rx_fifo/buff[73][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9821.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9822 (.I0(\i16/rx_fifo/buff[72][0] ), .I1(\i16/rx_fifo/buff[74][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9822.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9823 (.I0(n6155), .I1(n6156), .I2(n6122), .O(n6157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9823.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9824 (.I0(n6153), .I1(n6154), .I2(n6122), .I3(n6157), 
            .O(n6158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9824.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9825 (.I0(n6158), .I1(n6152), .I2(n6117), .I3(n6123), 
            .O(n6159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9825.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9826 (.I0(\i16/rx_fifo/buff[99][0] ), .I1(\i16/rx_fifo/buff[97][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9826.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9827 (.I0(\i16/rx_fifo/buff[96][0] ), .I1(\i16/rx_fifo/buff[98][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9827.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9828 (.I0(\i16/rx_fifo/buff[103][0] ), .I1(\i16/rx_fifo/buff[101][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9828.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9829 (.I0(\i16/rx_fifo/buff[100][0] ), .I1(\i16/rx_fifo/buff[102][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9829.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9830 (.I0(n6162), .I1(n6163), .I2(n6122), .I3(n6123), 
            .O(n6164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9830.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9831 (.I0(n6161), .I1(n6122), .I2(n6160), .I3(n6164), 
            .O(n6165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9831.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9832 (.I0(\i16/rx_fifo/buff[111][0] ), .I1(\i16/rx_fifo/buff[109][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9832.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9833 (.I0(\i16/rx_fifo/buff[108][0] ), .I1(\i16/rx_fifo/buff[110][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9833.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9834 (.I0(\i16/rx_fifo/buff[107][0] ), .I1(\i16/rx_fifo/buff[105][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9834.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9835 (.I0(\i16/rx_fifo/buff[104][0] ), .I1(\i16/rx_fifo/buff[106][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9835.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9836 (.I0(n6169), .I1(n6122), .I2(n6168), .I3(n6123), 
            .O(n6170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9836.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9837 (.I0(n6166), .I1(n6167), .I2(n6122), .I3(n6170), 
            .O(n6171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9837.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9838 (.I0(n6171), .I1(n6165), .I2(n6117), .I3(n6127), 
            .O(n6172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__9838.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__9839 (.I0(\i16/rx_fifo/buff[83][0] ), .I1(\i16/rx_fifo/buff[81][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9839.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9840 (.I0(\i16/rx_fifo/buff[80][0] ), .I1(\i16/rx_fifo/buff[82][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9840.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9841 (.I0(\i16/rx_fifo/buff[84][0] ), .I1(\i16/rx_fifo/buff[86][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9841.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9842 (.I0(n6173), .I1(n6174), .I2(n6175), .I3(n6122), 
            .O(n6176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__9842.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__9843 (.I0(\i16/rx_fifo/buff[87][0] ), .I1(\i16/rx_fifo/buff[85][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9843.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9844 (.I0(n6177), .I1(n6122), .I2(n6123), .I3(n6176), 
            .O(n6178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0c */ ;
    defparam LUT__9844.LUTMASK = 16'h0b0c;
    EFX_LUT4 LUT__9845 (.I0(\i16/rx_fifo/buff[91][0] ), .I1(\i16/rx_fifo/buff[89][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9845.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9846 (.I0(\i16/rx_fifo/buff[88][0] ), .I1(\i16/rx_fifo/buff[90][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9846.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9847 (.I0(\i16/rx_fifo/buff[95][0] ), .I1(\i16/rx_fifo/buff[93][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9847.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9848 (.I0(\i16/rx_fifo/buff[92][0] ), .I1(\i16/rx_fifo/buff[94][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9848.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9849 (.I0(n6181), .I1(n6182), .I2(n6122), .I3(n6123), 
            .O(n6183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9849.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9850 (.I0(n6180), .I1(n6122), .I2(n6179), .I3(n6183), 
            .O(n6184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9850.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9851 (.I0(n6114), .I1(n6118), .I2(ceg_net322), .O(n6185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__9851.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__9852 (.I0(n6178), .I1(n6184), .I2(n6117), .I3(n6185), 
            .O(n6186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9852.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9853 (.I0(\i16/rx_fifo/buff[127][0] ), .I1(\i16/rx_fifo/buff[125][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9853.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9854 (.I0(\i16/rx_fifo/buff[124][0] ), .I1(\i16/rx_fifo/buff[126][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9854.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9855 (.I0(\i16/rx_fifo/buff[123][0] ), .I1(\i16/rx_fifo/buff[121][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9855.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9856 (.I0(\i16/rx_fifo/buff[120][0] ), .I1(\i16/rx_fifo/buff[122][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9856.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9857 (.I0(n6189), .I1(n6190), .I2(n6188), .I3(n6122), 
            .O(n6191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__9857.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__9858 (.I0(n6187), .I1(n6122), .I2(n6191), .I3(n6123), 
            .O(n6192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__9858.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__9859 (.I0(\i16/rx_fifo/buff[116][0] ), .I1(\i16/rx_fifo/buff[118][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9859.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9860 (.I0(\i16/rx_fifo/buff[119][0] ), .I1(\i16/rx_fifo/buff[117][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6193), .O(n6194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9860.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9861 (.I0(\i16/rx_fifo/buff[115][0] ), .I1(\i16/rx_fifo/buff[113][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9861.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9862 (.I0(\i16/rx_fifo/buff[112][0] ), .I1(\i16/rx_fifo/buff[114][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9862.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9863 (.I0(n6196), .I1(n6122), .I2(n6195), .I3(n6123), 
            .O(n6197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9863.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9864 (.I0(n6194), .I1(n6122), .I2(n6197), .I3(n6117), 
            .O(n6198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__9864.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__9865 (.I0(n6192), .I1(n6198), .I2(n6127), .I3(n6185), 
            .O(n6199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__9865.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__9866 (.I0(n6186), .I1(n6199), .I2(n6159), .I3(n6172), 
            .O(n6200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__9866.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__9867 (.I0(rx_en_rx_packet), .I1(n6109), .O(n6201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9867.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9868 (.I0(\i16/rx_fifo/buff[55][0] ), .I1(\i16/rx_fifo/buff[53][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9868.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9869 (.I0(\i16/rx_fifo/buff[52][0] ), .I1(\i16/rx_fifo/buff[54][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9869.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9870 (.I0(\i16/rx_fifo/buff[51][0] ), .I1(\i16/rx_fifo/buff[49][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9870.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9871 (.I0(\i16/rx_fifo/buff[48][0] ), .I1(\i16/rx_fifo/buff[50][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9871.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9872 (.I0(n6205), .I1(n6122), .I2(n6204), .I3(n6123), 
            .O(n6206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9872.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9873 (.I0(n6202), .I1(n6203), .I2(n6122), .I3(n6206), 
            .O(n6207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9873.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9874 (.I0(\i16/rx_fifo/buff[60][0] ), .I1(\i16/rx_fifo/buff[62][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9874.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9875 (.I0(\i16/rx_fifo/buff[63][0] ), .I1(\i16/rx_fifo/buff[61][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6208), .O(n6209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9875.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9876 (.I0(\i16/rx_fifo/buff[59][0] ), .I1(\i16/rx_fifo/buff[57][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9876.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9877 (.I0(\i16/rx_fifo/buff[56][0] ), .I1(\i16/rx_fifo/buff[58][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9877.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9878 (.I0(n6211), .I1(n6122), .I2(n6210), .I3(n6123), 
            .O(n6212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9878.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9879 (.I0(n6209), .I1(n6122), .I2(n6212), .I3(n6127), 
            .O(n6213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__9879.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__9880 (.I0(\i16/rx_fifo/buff[39][0] ), .I1(\i16/rx_fifo/buff[37][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9880.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9881 (.I0(\i16/rx_fifo/buff[36][0] ), .I1(\i16/rx_fifo/buff[38][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9881.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9882 (.I0(\i16/rx_fifo/buff[35][0] ), .I1(\i16/rx_fifo/buff[33][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9882.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9883 (.I0(\i16/rx_fifo/buff[32][0] ), .I1(\i16/rx_fifo/buff[34][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9883.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9884 (.I0(n6217), .I1(n6122), .I2(n6216), .I3(n6123), 
            .O(n6218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9884.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9885 (.I0(n6214), .I1(n6215), .I2(n6122), .I3(n6218), 
            .O(n6219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9885.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9886 (.I0(\i16/rx_fifo/buff[44][0] ), .I1(\i16/rx_fifo/buff[46][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9886.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9887 (.I0(\i16/rx_fifo/buff[47][0] ), .I1(\i16/rx_fifo/buff[45][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6220), .O(n6221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9887.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9888 (.I0(\i16/rx_fifo/buff[43][0] ), .I1(\i16/rx_fifo/buff[41][0] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9888.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9889 (.I0(\i16/rx_fifo/buff[40][0] ), .I1(\i16/rx_fifo/buff[42][0] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9889.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9890 (.I0(n6223), .I1(n6122), .I2(n6222), .I3(n6123), 
            .O(n6224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9890.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9891 (.I0(n6221), .I1(n6122), .I2(n6224), .I3(n6127), 
            .O(n6225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__9891.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__9892 (.I0(n6219), .I1(n6225), .I2(n6207), .I3(n6213), 
            .O(n6226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__9892.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__9893 (.I0(n6114), .I1(n6118), .I2(ceg_net322), .I3(n6117), 
            .O(n6227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__9893.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__9894 (.I0(n6226), .I1(n6227), .I2(n6201), .I3(\rx_d[0] ), 
            .O(n6228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__9894.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__9895 (.I0(n6147), .I1(n6119), .I2(n6200), .I3(n6228), 
            .O(\rx_fifo/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4ff */ ;
    defparam LUT__9895.LUTMASK = 16'hf4ff;
    EFX_LUT4 LUT__9896 (.I0(n6114), .I1(n6109), .I2(rx_en_rx_packet_len), 
            .I3(n6115), .O(ceg_net498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__9896.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__9897 (.I0(rx_en_rx_packet_len), .I1(n193), .O(\rx_fifo/n152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__9897.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9898 (.I0(rx_en_rx_packet_len), .I1(n3196), .O(\rx_fifo/n151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__9898.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9899 (.I0(rx_en_rx_packet_len), .I1(n3192), .O(\rx_fifo/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__9899.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9900 (.I0(rx_en_rx_packet_len), .I1(n3189), .O(\rx_fifo/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__9900.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9901 (.I0(rx_en_rx_packet_len), .I1(n3185), .O(\rx_fifo/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__9901.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9902 (.I0(rx_en_rx_packet_len), .I1(n3182), .O(\rx_fifo/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__9902.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9903 (.I0(rx_en_rx_packet_len), .I1(n3179), .O(\rx_fifo/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__9903.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9904 (.I0(rx_en_rx_packet_len), .I1(\rx_fifo/rd_index[0] ), 
            .I2(\rx_fifo/rd_index[1] ), .O(\rx_fifo/n161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__9904.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__9905 (.I0(rx_en_rx_packet_len), .I1(n6122), .O(\rx_fifo/n160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__9905.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9906 (.I0(rx_en_rx_packet_len), .I1(n6123), .O(\rx_fifo/n159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__9906.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9907 (.I0(rx_en_rx_packet_len), .I1(n6127), .O(\rx_fifo/n158 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__9907.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9908 (.I0(rx_en_rx_packet_len), .I1(n6117), .O(\rx_fifo/n157 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__9908.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9909 (.I0(rx_en_rx_packet_len), .I1(n6118), .O(\rx_fifo/n156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__9909.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__9910 (.I0(n6118), .I1(\rx_fifo/rd_index[6] ), .I2(rx_en_rx_packet_len), 
            .I3(\rx_fifo/rd_index[7] ), .O(\rx_fifo/n155 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b04 */ ;
    defparam LUT__9910.LUTMASK = 16'h0b04;
    EFX_LUT4 LUT__9911 (.I0(rx_en_rx_packet_len), .I1(\rx_d[1] ), .O(\data_to_rx_packet_len_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9911.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9912 (.I0(rx_en_rx_packet_len), .I1(\rx_d[2] ), .O(\data_to_rx_packet_len_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9912.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9913 (.I0(rx_en_rx_packet_len), .I1(\rx_d[3] ), .O(\data_to_rx_packet_len_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9913.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9914 (.I0(rx_en_rx_packet_len), .I1(\rx_d[4] ), .O(\data_to_rx_packet_len_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9914.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9915 (.I0(rx_en_rx_packet_len), .I1(\rx_d[5] ), .O(\data_to_rx_packet_len_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9915.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9916 (.I0(rx_en_rx_packet_len), .I1(\rx_d[6] ), .O(\data_to_rx_packet_len_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9916.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9917 (.I0(rx_en_rx_packet_len), .I1(\rx_d[7] ), .O(\data_to_rx_packet_len_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__9917.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__9918 (.I0(\i16/rx_fifo/buff[7][1] ), .I1(\i16/rx_fifo/buff[5][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9918.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9919 (.I0(\i16/rx_fifo/buff[4][1] ), .I1(\i16/rx_fifo/buff[6][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9919.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9920 (.I0(n6229), .I1(n6230), .I2(n6122), .O(n6231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__9920.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__9921 (.I0(\i16/rx_fifo/buff[3][1] ), .I1(\i16/rx_fifo/buff[1][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9921.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9922 (.I0(\i16/rx_fifo/buff[0][1] ), .I1(\i16/rx_fifo/buff[2][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9922.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9923 (.I0(n6233), .I1(n6122), .I2(n6232), .I3(n6123), 
            .O(n6234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9923.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9924 (.I0(\i16/rx_fifo/buff[11][1] ), .I1(\i16/rx_fifo/buff[9][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9924.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9925 (.I0(\i16/rx_fifo/buff[8][1] ), .I1(\i16/rx_fifo/buff[10][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9925.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9926 (.I0(n6235), .I1(n6236), .I2(n6122), .O(n6237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__9926.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__9927 (.I0(\i16/rx_fifo/buff[15][1] ), .I1(\i16/rx_fifo/buff[13][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9927.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9928 (.I0(\i16/rx_fifo/buff[12][1] ), .I1(\i16/rx_fifo/buff[14][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9928.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9929 (.I0(n6238), .I1(n6239), .I2(n6122), .I3(n6123), 
            .O(n6240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9929.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9930 (.I0(n6237), .I1(n6240), .I2(n6231), .I3(n6234), 
            .O(n6241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__9930.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__9931 (.I0(\i16/rx_fifo/buff[39][1] ), .I1(\i16/rx_fifo/buff[37][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9931.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9932 (.I0(\i16/rx_fifo/buff[36][1] ), .I1(\i16/rx_fifo/buff[38][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9932.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9933 (.I0(n6242), .I1(n6243), .I2(n6122), .O(n6244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__9933.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__9934 (.I0(\i16/rx_fifo/buff[35][1] ), .I1(\i16/rx_fifo/buff[33][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9934.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9935 (.I0(\i16/rx_fifo/buff[32][1] ), .I1(\i16/rx_fifo/buff[34][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9935.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9936 (.I0(n6246), .I1(n6122), .I2(n6245), .I3(n6123), 
            .O(n6247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9936.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9937 (.I0(\i16/rx_fifo/buff[47][1] ), .I1(\i16/rx_fifo/buff[45][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9937.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9938 (.I0(\i16/rx_fifo/buff[44][1] ), .I1(\i16/rx_fifo/buff[46][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9938.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9939 (.I0(n6248), .I1(n6249), .I2(n6122), .O(n6250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__9939.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__9940 (.I0(\i16/rx_fifo/buff[43][1] ), .I1(\i16/rx_fifo/buff[41][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9940.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9941 (.I0(\i16/rx_fifo/buff[40][1] ), .I1(\i16/rx_fifo/buff[42][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9941.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9942 (.I0(n6252), .I1(n6122), .I2(n6251), .I3(n6123), 
            .O(n6253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9942.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9943 (.I0(n6250), .I1(n6253), .I2(n6244), .I3(n6247), 
            .O(n6254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__9943.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__9944 (.I0(n6254), .I1(n6241), .I2(n6127), .I3(n6117), 
            .O(n6255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9944.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9945 (.I0(n6255), .I1(n6114), .I2(n6118), .I3(ceg_net322), 
            .O(n6256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__9945.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__9946 (.I0(\i16/rx_fifo/buff[20][1] ), .I1(\i16/rx_fifo/buff[22][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9946.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9947 (.I0(\i16/rx_fifo/buff[23][1] ), .I1(\i16/rx_fifo/buff[21][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6257), .O(n6258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9947.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9948 (.I0(\i16/rx_fifo/buff[16][1] ), .I1(\i16/rx_fifo/buff[18][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__9948.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__9949 (.I0(\i16/rx_fifo/buff[19][1] ), .I1(\i16/rx_fifo/buff[17][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6259), .O(n6260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__9949.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__9950 (.I0(n6260), .I1(n6258), .I2(n6123), .I3(n6122), 
            .O(n6261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__9950.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__9951 (.I0(\i16/rx_fifo/buff[55][1] ), .I1(\i16/rx_fifo/buff[53][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9951.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9952 (.I0(\i16/rx_fifo/buff[52][1] ), .I1(\i16/rx_fifo/buff[54][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9952.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9953 (.I0(\i16/rx_fifo/buff[51][1] ), .I1(\i16/rx_fifo/buff[49][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9953.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9954 (.I0(\i16/rx_fifo/buff[48][1] ), .I1(\i16/rx_fifo/buff[50][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9954.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9955 (.I0(n6265), .I1(n6122), .I2(n6264), .I3(n6123), 
            .O(n6266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9955.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9956 (.I0(n6262), .I1(n6263), .I2(n6122), .I3(n6266), 
            .O(n6267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9956.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9957 (.I0(\i16/rx_fifo/buff[63][1] ), .I1(\i16/rx_fifo/buff[61][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9957.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9958 (.I0(\i16/rx_fifo/buff[60][1] ), .I1(\i16/rx_fifo/buff[62][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9958.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9959 (.I0(\i16/rx_fifo/buff[59][1] ), .I1(\i16/rx_fifo/buff[57][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9959.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9960 (.I0(\i16/rx_fifo/buff[56][1] ), .I1(\i16/rx_fifo/buff[58][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9960.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9961 (.I0(n6271), .I1(n6122), .I2(n6270), .I3(n6123), 
            .O(n6272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9961.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9962 (.I0(n6268), .I1(n6269), .I2(n6122), .I3(n6272), 
            .O(n6273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9962.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9963 (.I0(n6273), .I1(n6267), .I2(\rx_fifo/rd_index[5] ), 
            .I3(n6127), .O(n6274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9963.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9964 (.I0(\i16/rx_fifo/buff[31][1] ), .I1(\i16/rx_fifo/buff[29][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9964.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9965 (.I0(\i16/rx_fifo/buff[28][1] ), .I1(\i16/rx_fifo/buff[30][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9965.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9966 (.I0(\i16/rx_fifo/buff[27][1] ), .I1(\i16/rx_fifo/buff[25][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9966.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9967 (.I0(\i16/rx_fifo/buff[24][1] ), .I1(\i16/rx_fifo/buff[26][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9967.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9968 (.I0(n6278), .I1(n6122), .I2(n6277), .I3(n6123), 
            .O(n6279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9968.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9969 (.I0(n6275), .I1(n6276), .I2(n6122), .I3(n6279), 
            .O(n6280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__9969.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__9970 (.I0(\rx_fifo/rd_index[5] ), .I1(n6261), .I2(n6280), 
            .I3(n6274), .O(n6281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__9970.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__9971 (.I0(\i16/rx_fifo/buff[92][1] ), .I1(\i16/rx_fifo/buff[94][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9971.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9972 (.I0(\i16/rx_fifo/buff[91][1] ), .I1(\i16/rx_fifo/buff[89][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9972.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9973 (.I0(\i16/rx_fifo/buff[88][1] ), .I1(\i16/rx_fifo/buff[90][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9973.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9974 (.I0(n6283), .I1(n6284), .I2(n6282), .I3(n6122), 
            .O(n6285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__9974.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__9975 (.I0(n6285), .I1(n6123), .I2(n6127), .O(n6286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__9975.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__9976 (.I0(\i16/rx_fifo/buff[83][1] ), .I1(\i16/rx_fifo/buff[81][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9976.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9977 (.I0(\i16/rx_fifo/buff[80][1] ), .I1(\i16/rx_fifo/buff[82][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9977.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9978 (.I0(\i16/rx_fifo/buff[87][1] ), .I1(\i16/rx_fifo/buff[85][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9978.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9979 (.I0(\i16/rx_fifo/buff[84][1] ), .I1(\i16/rx_fifo/buff[86][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9979.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9980 (.I0(\i16/rx_fifo/buff[95][1] ), .I1(\i16/rx_fifo/buff[93][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9980.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9981 (.I0(n6289), .I1(n6290), .I2(n6291), .I3(n6123), 
            .O(n6292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__9981.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__9982 (.I0(n6287), .I1(n6288), .I2(n6292), .I3(n6122), 
            .O(n6293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__9982.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__9983 (.I0(n6122), .I1(n6123), .I2(n6293), .I3(n6286), 
            .O(n6294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc700 */ ;
    defparam LUT__9983.LUTMASK = 16'hc700;
    EFX_LUT4 LUT__9984 (.I0(\i16/rx_fifo/buff[79][1] ), .I1(\i16/rx_fifo/buff[77][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9984.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9985 (.I0(\i16/rx_fifo/buff[76][1] ), .I1(\i16/rx_fifo/buff[78][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9985.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9986 (.I0(\i16/rx_fifo/buff[75][1] ), .I1(\i16/rx_fifo/buff[73][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9986.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9987 (.I0(\i16/rx_fifo/buff[72][1] ), .I1(\i16/rx_fifo/buff[74][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9987.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9988 (.I0(n6297), .I1(n6298), .I2(n6296), .I3(n6122), 
            .O(n6299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__9988.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__9989 (.I0(n6295), .I1(n6122), .I2(n6299), .I3(n6123), 
            .O(n6300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__9989.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__9990 (.I0(\i16/rx_fifo/buff[71][1] ), .I1(\i16/rx_fifo/buff[69][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9990.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9991 (.I0(\i16/rx_fifo/buff[68][1] ), .I1(\i16/rx_fifo/buff[70][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9991.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9992 (.I0(\i16/rx_fifo/buff[67][1] ), .I1(\i16/rx_fifo/buff[65][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9992.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9993 (.I0(\i16/rx_fifo/buff[64][1] ), .I1(\i16/rx_fifo/buff[66][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9993.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9994 (.I0(n6303), .I1(n6304), .I2(n6302), .I3(n6122), 
            .O(n6305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__9994.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__9995 (.I0(n6301), .I1(n6122), .I2(n6123), .I3(n6305), 
            .O(n6306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0c */ ;
    defparam LUT__9995.LUTMASK = 16'h0b0c;
    EFX_LUT4 LUT__9996 (.I0(n6300), .I1(n6127), .I2(n6306), .I3(n6117), 
            .O(n6307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__9996.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__9997 (.I0(\i16/rx_fifo/buff[107][1] ), .I1(\i16/rx_fifo/buff[105][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__9997.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__9998 (.I0(\i16/rx_fifo/buff[104][1] ), .I1(\i16/rx_fifo/buff[106][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9998.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__9999 (.I0(\i16/rx_fifo/buff[108][1] ), .I1(\i16/rx_fifo/buff[110][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__9999.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10000 (.I0(n6308), .I1(n6309), .I2(n6310), .I3(n6122), 
            .O(n6311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10000.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10001 (.I0(\i16/rx_fifo/buff[111][1] ), .I1(\i16/rx_fifo/buff[109][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10001.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10002 (.I0(n6312), .I1(n6122), .I2(n6311), .I3(n6123), 
            .O(n6313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__10002.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__10003 (.I0(\i16/rx_fifo/buff[103][1] ), .I1(\i16/rx_fifo/buff[101][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10003.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10004 (.I0(\i16/rx_fifo/buff[100][1] ), .I1(\i16/rx_fifo/buff[102][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10004.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10005 (.I0(\i16/rx_fifo/buff[99][1] ), .I1(\i16/rx_fifo/buff[97][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10005.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10006 (.I0(\i16/rx_fifo/buff[96][1] ), .I1(\i16/rx_fifo/buff[98][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10006.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10007 (.I0(n6316), .I1(n6317), .I2(n6315), .I3(n6122), 
            .O(n6318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10007.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10008 (.I0(n6314), .I1(n6122), .I2(n6123), .I3(n6318), 
            .O(n6319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0c */ ;
    defparam LUT__10008.LUTMASK = 16'h0b0c;
    EFX_LUT4 LUT__10009 (.I0(n6313), .I1(n6127), .I2(n6319), .I3(n6185), 
            .O(n6320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10009.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10010 (.I0(\i16/rx_fifo/buff[127][1] ), .I1(\i16/rx_fifo/buff[125][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10010.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10011 (.I0(\i16/rx_fifo/buff[124][1] ), .I1(\i16/rx_fifo/buff[126][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10011.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10012 (.I0(n6321), .I1(n6322), .I2(n6122), .O(n6323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10012.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10013 (.I0(\i16/rx_fifo/buff[123][1] ), .I1(\i16/rx_fifo/buff[121][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10013.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10014 (.I0(\i16/rx_fifo/buff[120][1] ), .I1(\i16/rx_fifo/buff[122][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10014.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10015 (.I0(n6325), .I1(n6122), .I2(n6324), .I3(n6123), 
            .O(n6326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10015.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10016 (.I0(\i16/rx_fifo/buff[119][1] ), .I1(\i16/rx_fifo/buff[117][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10016.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10017 (.I0(\i16/rx_fifo/buff[116][1] ), .I1(\i16/rx_fifo/buff[118][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10017.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10018 (.I0(n6327), .I1(n6328), .I2(n6122), .O(n6329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10018.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10019 (.I0(\i16/rx_fifo/buff[115][1] ), .I1(\i16/rx_fifo/buff[113][1] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10019.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10020 (.I0(\i16/rx_fifo/buff[112][1] ), .I1(\i16/rx_fifo/buff[114][1] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10020.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10021 (.I0(n6331), .I1(n6122), .I2(n6330), .I3(n6123), 
            .O(n6332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10021.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10022 (.I0(n6329), .I1(n6332), .I2(n6323), .I3(n6326), 
            .O(n6333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10022.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10023 (.I0(n6333), .I1(n6127), .I2(n6117), .I3(n6185), 
            .O(n6334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__10023.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__10024 (.I0(n6320), .I1(n6334), .I2(n6294), .I3(n6307), 
            .O(n6335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__10024.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__10025 (.I0(n6201), .I1(\rx_d[1] ), .O(n6336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10025.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10026 (.I0(n6281), .I1(n6256), .I2(n6335), .I3(n6336), 
            .O(\rx_fifo/n143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4 */ ;
    defparam LUT__10026.LUTMASK = 16'hfff4;
    EFX_LUT4 LUT__10027 (.I0(\i16/rx_fifo/buff[79][2] ), .I1(\i16/rx_fifo/buff[77][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10027.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10028 (.I0(\i16/rx_fifo/buff[76][2] ), .I1(\i16/rx_fifo/buff[78][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10028.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10029 (.I0(n6337), .I1(n6338), .I2(n6122), .O(n6339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10029.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10030 (.I0(\i16/rx_fifo/buff[75][2] ), .I1(\i16/rx_fifo/buff[73][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10030.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10031 (.I0(\i16/rx_fifo/buff[72][2] ), .I1(\i16/rx_fifo/buff[74][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10031.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10032 (.I0(n6341), .I1(n6122), .I2(n6340), .I3(n6123), 
            .O(n6342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10032.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10033 (.I0(\i16/rx_fifo/buff[71][2] ), .I1(\i16/rx_fifo/buff[69][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10033.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10034 (.I0(\i16/rx_fifo/buff[68][2] ), .I1(\i16/rx_fifo/buff[70][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10034.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10035 (.I0(n6343), .I1(n6344), .I2(n6122), .O(n6345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10035.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10036 (.I0(\i16/rx_fifo/buff[67][2] ), .I1(\i16/rx_fifo/buff[65][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10036.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10037 (.I0(\i16/rx_fifo/buff[64][2] ), .I1(\i16/rx_fifo/buff[66][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10037.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10038 (.I0(n6347), .I1(n6122), .I2(n6346), .I3(n6123), 
            .O(n6348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10038.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10039 (.I0(n6345), .I1(n6348), .I2(n6339), .I3(n6342), 
            .O(n6349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10039.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10040 (.I0(\i16/rx_fifo/buff[111][2] ), .I1(\i16/rx_fifo/buff[109][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10040.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10041 (.I0(\i16/rx_fifo/buff[108][2] ), .I1(\i16/rx_fifo/buff[110][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10041.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10042 (.I0(n6350), .I1(n6351), .I2(n6122), .O(n6352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10042.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10043 (.I0(\i16/rx_fifo/buff[107][2] ), .I1(\i16/rx_fifo/buff[105][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10043.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10044 (.I0(\i16/rx_fifo/buff[104][2] ), .I1(\i16/rx_fifo/buff[106][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10044.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10045 (.I0(n6354), .I1(n6122), .I2(n6353), .I3(n6123), 
            .O(n6355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10045.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10046 (.I0(\i16/rx_fifo/buff[103][2] ), .I1(\i16/rx_fifo/buff[101][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10046.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10047 (.I0(\i16/rx_fifo/buff[100][2] ), .I1(\i16/rx_fifo/buff[102][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10047.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10048 (.I0(n6356), .I1(n6357), .I2(n6122), .O(n6358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10048.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10049 (.I0(\i16/rx_fifo/buff[99][2] ), .I1(\i16/rx_fifo/buff[97][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10049.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10050 (.I0(\i16/rx_fifo/buff[96][2] ), .I1(\i16/rx_fifo/buff[98][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10050.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10051 (.I0(n6360), .I1(n6122), .I2(n6359), .I3(n6123), 
            .O(n6361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10051.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10052 (.I0(n6358), .I1(n6361), .I2(n6352), .I3(n6355), 
            .O(n6362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10052.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10053 (.I0(n6362), .I1(n6349), .I2(n6127), .I3(n6117), 
            .O(n6363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10053.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10054 (.I0(\i16/rx_fifo/buff[83][2] ), .I1(\i16/rx_fifo/buff[81][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10054.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10055 (.I0(\i16/rx_fifo/buff[80][2] ), .I1(\i16/rx_fifo/buff[82][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10055.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10056 (.I0(n6364), .I1(n6365), .I2(n6122), .O(n6366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10056.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10057 (.I0(\i16/rx_fifo/buff[87][2] ), .I1(\i16/rx_fifo/buff[85][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10057.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10058 (.I0(\i16/rx_fifo/buff[84][2] ), .I1(\i16/rx_fifo/buff[86][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10058.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10059 (.I0(n6367), .I1(n6368), .I2(n6122), .I3(n6123), 
            .O(n6369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10059.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10060 (.I0(\i16/rx_fifo/buff[95][2] ), .I1(\i16/rx_fifo/buff[93][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10060.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10061 (.I0(\i16/rx_fifo/buff[92][2] ), .I1(\i16/rx_fifo/buff[94][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10061.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10062 (.I0(n6370), .I1(n6371), .I2(n6122), .O(n6372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10062.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10063 (.I0(\i16/rx_fifo/buff[91][2] ), .I1(\i16/rx_fifo/buff[89][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10063.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10064 (.I0(\i16/rx_fifo/buff[88][2] ), .I1(\i16/rx_fifo/buff[90][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10064.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10065 (.I0(n6374), .I1(n6122), .I2(n6373), .I3(n6123), 
            .O(n6375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10065.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10066 (.I0(n6372), .I1(n6375), .I2(n6366), .I3(n6369), 
            .O(n6376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10066.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10067 (.I0(\i16/rx_fifo/buff[127][2] ), .I1(\i16/rx_fifo/buff[125][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10067.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10068 (.I0(\i16/rx_fifo/buff[124][2] ), .I1(\i16/rx_fifo/buff[126][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10068.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10069 (.I0(n6377), .I1(n6378), .I2(n6122), .O(n6379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10069.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10070 (.I0(\i16/rx_fifo/buff[123][2] ), .I1(\i16/rx_fifo/buff[121][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10070.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10071 (.I0(\i16/rx_fifo/buff[120][2] ), .I1(\i16/rx_fifo/buff[122][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10071.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10072 (.I0(n6381), .I1(n6122), .I2(n6380), .I3(n6123), 
            .O(n6382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10072.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10073 (.I0(\i16/rx_fifo/buff[119][2] ), .I1(\i16/rx_fifo/buff[117][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10073.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10074 (.I0(\i16/rx_fifo/buff[116][2] ), .I1(\i16/rx_fifo/buff[118][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10074.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10075 (.I0(n6383), .I1(n6384), .I2(n6122), .O(n6385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10075.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10076 (.I0(\i16/rx_fifo/buff[115][2] ), .I1(\i16/rx_fifo/buff[113][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10076.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10077 (.I0(\i16/rx_fifo/buff[112][2] ), .I1(\i16/rx_fifo/buff[114][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10077.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10078 (.I0(n6387), .I1(n6122), .I2(n6386), .I3(n6123), 
            .O(n6388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10078.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10079 (.I0(n6385), .I1(n6388), .I2(n6379), .I3(n6382), 
            .O(n6389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10079.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10080 (.I0(n6389), .I1(n6376), .I2(\rx_fifo/rd_index[5] ), 
            .I3(n6127), .O(n6390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10080.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10081 (.I0(n6363), .I1(n6390), .I2(n6185), .O(n6391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10081.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10082 (.I0(\i16/rx_fifo/buff[39][2] ), .I1(\i16/rx_fifo/buff[37][2] ), 
            .I2(n6123), .I3(\rx_fifo/rd_index[1] ), .O(n6392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__10082.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__10083 (.I0(\i16/rx_fifo/buff[47][2] ), .I1(\i16/rx_fifo/buff[45][2] ), 
            .I2(n6123), .I3(n6392), .O(n6393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcfa0 */ ;
    defparam LUT__10083.LUTMASK = 16'hcfa0;
    EFX_LUT4 LUT__10084 (.I0(\i16/rx_fifo/buff[36][2] ), .I1(\i16/rx_fifo/buff[38][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10084.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10085 (.I0(\i16/rx_fifo/buff[35][2] ), .I1(\i16/rx_fifo/buff[33][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10085.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10086 (.I0(\i16/rx_fifo/buff[32][2] ), .I1(\i16/rx_fifo/buff[34][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10086.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10087 (.I0(n6395), .I1(n6396), .I2(n6394), .I3(n6122), 
            .O(n6397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10087.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10088 (.I0(\i16/rx_fifo/buff[43][2] ), .I1(\i16/rx_fifo/buff[41][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10088.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10089 (.I0(\i16/rx_fifo/buff[40][2] ), .I1(\i16/rx_fifo/buff[42][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10089.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10090 (.I0(\i16/rx_fifo/buff[44][2] ), .I1(\i16/rx_fifo/buff[46][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10090.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10091 (.I0(n6398), .I1(n6399), .I2(n6400), .I3(n6122), 
            .O(n6401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10091.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10092 (.I0(n6397), .I1(n6401), .I2(n6123), .O(n6402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__10092.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__10093 (.I0(n6393), .I1(\rx_fifo/rd_index[0] ), .I2(n6402), 
            .I3(n6122), .O(n6403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ef0 */ ;
    defparam LUT__10093.LUTMASK = 16'h0ef0;
    EFX_LUT4 LUT__10094 (.I0(n6114), .I1(n6118), .I2(n6127), .I3(ceg_net322), 
            .O(n6404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10094.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10095 (.I0(n6114), .I1(n6118), .I2(n6127), .I3(ceg_net322), 
            .O(n6405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10095.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10096 (.I0(\i16/rx_fifo/buff[51][2] ), .I1(\i16/rx_fifo/buff[49][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10096.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10097 (.I0(\i16/rx_fifo/buff[48][2] ), .I1(\i16/rx_fifo/buff[50][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10097.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10098 (.I0(n6406), .I1(n6407), .I2(n6122), .O(n6408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10098.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10099 (.I0(\i16/rx_fifo/buff[55][2] ), .I1(\i16/rx_fifo/buff[53][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10099.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10100 (.I0(\i16/rx_fifo/buff[52][2] ), .I1(\i16/rx_fifo/buff[54][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10100.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10101 (.I0(n6409), .I1(n6410), .I2(n6122), .I3(n6123), 
            .O(n6411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10101.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10102 (.I0(\i16/rx_fifo/buff[63][2] ), .I1(\i16/rx_fifo/buff[61][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10102.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10103 (.I0(\i16/rx_fifo/buff[60][2] ), .I1(\i16/rx_fifo/buff[62][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10103.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10104 (.I0(n6412), .I1(n6413), .I2(n6122), .O(n6414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10104.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10105 (.I0(\i16/rx_fifo/buff[59][2] ), .I1(\i16/rx_fifo/buff[57][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10105.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10106 (.I0(\i16/rx_fifo/buff[56][2] ), .I1(\i16/rx_fifo/buff[58][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10106.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10107 (.I0(n6416), .I1(n6122), .I2(n6415), .I3(n6123), 
            .O(n6417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10107.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10108 (.I0(n6414), .I1(n6417), .I2(n6408), .I3(n6411), 
            .O(n6418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10108.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10109 (.I0(n6418), .I1(n6405), .I2(n6119), .O(n6419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__10109.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__10110 (.I0(\i16/rx_fifo/buff[15][2] ), .I1(\i16/rx_fifo/buff[13][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10110.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10111 (.I0(\i16/rx_fifo/buff[12][2] ), .I1(\i16/rx_fifo/buff[14][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10111.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10112 (.I0(n6420), .I1(n6421), .I2(n6122), .O(n6422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10112.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10113 (.I0(\i16/rx_fifo/buff[11][2] ), .I1(\i16/rx_fifo/buff[9][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10113.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10114 (.I0(\i16/rx_fifo/buff[8][2] ), .I1(\i16/rx_fifo/buff[10][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10114.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10115 (.I0(n6424), .I1(n6122), .I2(n6423), .I3(n6123), 
            .O(n6425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10115.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10116 (.I0(\i16/rx_fifo/buff[7][2] ), .I1(\i16/rx_fifo/buff[5][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10116.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10117 (.I0(\i16/rx_fifo/buff[4][2] ), .I1(\i16/rx_fifo/buff[6][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10117.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10118 (.I0(n6426), .I1(n6427), .I2(n6122), .O(n6428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10118.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10119 (.I0(\i16/rx_fifo/buff[3][2] ), .I1(\i16/rx_fifo/buff[1][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10119.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10120 (.I0(\i16/rx_fifo/buff[0][2] ), .I1(\i16/rx_fifo/buff[2][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10120.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10121 (.I0(n6430), .I1(n6122), .I2(n6429), .I3(n6123), 
            .O(n6431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10121.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10122 (.I0(n6428), .I1(n6431), .I2(n6422), .I3(n6425), 
            .O(n6432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10122.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10123 (.I0(\i16/rx_fifo/buff[31][2] ), .I1(\i16/rx_fifo/buff[29][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10123.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10124 (.I0(\i16/rx_fifo/buff[28][2] ), .I1(\i16/rx_fifo/buff[30][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10124.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10125 (.I0(n6433), .I1(n6434), .I2(n6122), .O(n6435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10125.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10126 (.I0(\i16/rx_fifo/buff[27][2] ), .I1(\i16/rx_fifo/buff[25][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10126.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10127 (.I0(\i16/rx_fifo/buff[24][2] ), .I1(\i16/rx_fifo/buff[26][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10127.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10128 (.I0(n6437), .I1(n6122), .I2(n6436), .I3(n6123), 
            .O(n6438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10128.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10129 (.I0(\i16/rx_fifo/buff[23][2] ), .I1(\i16/rx_fifo/buff[21][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10129.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10130 (.I0(\i16/rx_fifo/buff[20][2] ), .I1(\i16/rx_fifo/buff[22][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10130.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10131 (.I0(n6439), .I1(n6440), .I2(n6122), .O(n6441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10131.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10132 (.I0(\i16/rx_fifo/buff[19][2] ), .I1(\i16/rx_fifo/buff[17][2] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10132.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10133 (.I0(\i16/rx_fifo/buff[16][2] ), .I1(\i16/rx_fifo/buff[18][2] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10133.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10134 (.I0(n6443), .I1(n6122), .I2(n6442), .I3(n6123), 
            .O(n6444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10134.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10135 (.I0(n6441), .I1(n6444), .I2(n6435), .I3(n6438), 
            .O(n6445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10135.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10136 (.I0(n6445), .I1(n6432), .I2(n6117), .I3(n6127), 
            .O(n6446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10136.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10137 (.I0(n6404), .I1(n6403), .I2(n6419), .I3(n6446), 
            .O(n6447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__10137.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__10138 (.I0(n6201), .I1(\rx_d[2] ), .I2(n6391), .I3(n6447), 
            .O(\rx_fifo/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__10138.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__10139 (.I0(\i16/rx_fifo/buff[71][3] ), .I1(\i16/rx_fifo/buff[69][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10139.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10140 (.I0(\i16/rx_fifo/buff[68][3] ), .I1(\i16/rx_fifo/buff[70][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10140.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10141 (.I0(n6448), .I1(n6449), .I2(n6122), .O(n6450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10141.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10142 (.I0(\i16/rx_fifo/buff[67][3] ), .I1(\i16/rx_fifo/buff[65][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10142.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10143 (.I0(\i16/rx_fifo/buff[64][3] ), .I1(\i16/rx_fifo/buff[66][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10143.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10144 (.I0(n6452), .I1(n6122), .I2(n6451), .I3(n6123), 
            .O(n6453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10144.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10145 (.I0(\i16/rx_fifo/buff[79][3] ), .I1(\i16/rx_fifo/buff[77][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10145.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10146 (.I0(\i16/rx_fifo/buff[76][3] ), .I1(\i16/rx_fifo/buff[78][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10146.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10147 (.I0(n6454), .I1(n6455), .I2(n6122), .O(n6456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10147.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10148 (.I0(\i16/rx_fifo/buff[75][3] ), .I1(\i16/rx_fifo/buff[73][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10148.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10149 (.I0(\i16/rx_fifo/buff[72][3] ), .I1(\i16/rx_fifo/buff[74][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10149.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10150 (.I0(n6458), .I1(n6122), .I2(n6457), .I3(n6123), 
            .O(n6459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10150.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10151 (.I0(n6456), .I1(n6459), .I2(n6450), .I3(n6453), 
            .O(n6460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10151.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10152 (.I0(\i16/rx_fifo/buff[111][3] ), .I1(\i16/rx_fifo/buff[109][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10152.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10153 (.I0(\i16/rx_fifo/buff[108][3] ), .I1(\i16/rx_fifo/buff[110][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10153.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10154 (.I0(n6461), .I1(n6462), .I2(n6122), .O(n6463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10154.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10155 (.I0(\i16/rx_fifo/buff[107][3] ), .I1(\i16/rx_fifo/buff[105][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10155.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10156 (.I0(\i16/rx_fifo/buff[104][3] ), .I1(\i16/rx_fifo/buff[106][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10156.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10157 (.I0(n6465), .I1(n6122), .I2(n6464), .I3(n6123), 
            .O(n6466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10157.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10158 (.I0(\i16/rx_fifo/buff[103][3] ), .I1(\i16/rx_fifo/buff[101][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10158.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10159 (.I0(\i16/rx_fifo/buff[100][3] ), .I1(\i16/rx_fifo/buff[102][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10159.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10160 (.I0(n6467), .I1(n6468), .I2(n6122), .O(n6469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10160.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10161 (.I0(\i16/rx_fifo/buff[99][3] ), .I1(\i16/rx_fifo/buff[97][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10161.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10162 (.I0(\i16/rx_fifo/buff[96][3] ), .I1(\i16/rx_fifo/buff[98][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10162.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10163 (.I0(n6471), .I1(n6122), .I2(n6470), .I3(n6123), 
            .O(n6472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10163.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10164 (.I0(n6469), .I1(n6472), .I2(n6463), .I3(n6466), 
            .O(n6473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10164.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10165 (.I0(n6473), .I1(n6460), .I2(n6127), .I3(n6117), 
            .O(n6474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10165.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10166 (.I0(\i16/rx_fifo/buff[119][3] ), .I1(\i16/rx_fifo/buff[117][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10166.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10167 (.I0(\i16/rx_fifo/buff[116][3] ), .I1(\i16/rx_fifo/buff[118][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10167.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10168 (.I0(n6475), .I1(n6476), .I2(n6122), .O(n6477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10168.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10169 (.I0(\i16/rx_fifo/buff[115][3] ), .I1(\i16/rx_fifo/buff[113][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10169.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10170 (.I0(\i16/rx_fifo/buff[112][3] ), .I1(\i16/rx_fifo/buff[114][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10170.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10171 (.I0(n6479), .I1(n6122), .I2(n6478), .I3(n6123), 
            .O(n6480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10171.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10172 (.I0(\i16/rx_fifo/buff[127][3] ), .I1(\i16/rx_fifo/buff[125][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10172.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10173 (.I0(\i16/rx_fifo/buff[124][3] ), .I1(\i16/rx_fifo/buff[126][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10173.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10174 (.I0(n6481), .I1(n6482), .I2(n6122), .O(n6483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10174.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10175 (.I0(\i16/rx_fifo/buff[123][3] ), .I1(\i16/rx_fifo/buff[121][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10175.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10176 (.I0(\i16/rx_fifo/buff[120][3] ), .I1(\i16/rx_fifo/buff[122][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10176.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10177 (.I0(n6485), .I1(n6122), .I2(n6484), .I3(n6123), 
            .O(n6486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10177.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10178 (.I0(n6483), .I1(n6486), .I2(n6477), .I3(n6480), 
            .O(n6487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10178.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10179 (.I0(\i16/rx_fifo/buff[83][3] ), .I1(\i16/rx_fifo/buff[81][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10179.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10180 (.I0(\i16/rx_fifo/buff[80][3] ), .I1(\i16/rx_fifo/buff[82][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10180.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10181 (.I0(n6488), .I1(n6489), .I2(n6122), .O(n6490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10181.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10182 (.I0(\i16/rx_fifo/buff[87][3] ), .I1(\i16/rx_fifo/buff[85][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10182.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10183 (.I0(\i16/rx_fifo/buff[84][3] ), .I1(\i16/rx_fifo/buff[86][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10183.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10184 (.I0(n6491), .I1(n6492), .I2(n6122), .I3(n6123), 
            .O(n6493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10184.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10185 (.I0(\i16/rx_fifo/buff[95][3] ), .I1(\i16/rx_fifo/buff[93][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10185.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10186 (.I0(\i16/rx_fifo/buff[92][3] ), .I1(\i16/rx_fifo/buff[94][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10186.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10187 (.I0(n6494), .I1(n6495), .I2(n6122), .O(n6496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10187.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10188 (.I0(\i16/rx_fifo/buff[91][3] ), .I1(\i16/rx_fifo/buff[89][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10188.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10189 (.I0(\i16/rx_fifo/buff[88][3] ), .I1(\i16/rx_fifo/buff[90][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10189.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10190 (.I0(n6498), .I1(n6122), .I2(n6497), .I3(n6123), 
            .O(n6499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10190.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10191 (.I0(n6496), .I1(n6499), .I2(n6490), .I3(n6493), 
            .O(n6500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10191.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10192 (.I0(n6500), .I1(n6487), .I2(\rx_fifo/rd_index[5] ), 
            .I3(n6127), .O(n6501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__10192.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__10193 (.I0(n6474), .I1(n6501), .I2(n6185), .O(n6502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10193.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10194 (.I0(\i16/rx_fifo/buff[31][3] ), .I1(\i16/rx_fifo/buff[29][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10194.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10195 (.I0(\i16/rx_fifo/buff[28][3] ), .I1(\i16/rx_fifo/buff[30][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10195.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10196 (.I0(\i16/rx_fifo/buff[27][3] ), .I1(\i16/rx_fifo/buff[25][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10196.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10197 (.I0(\i16/rx_fifo/buff[24][3] ), .I1(\i16/rx_fifo/buff[26][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10197.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10198 (.I0(n6505), .I1(n6506), .I2(n6504), .I3(n6122), 
            .O(n6507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10198.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10199 (.I0(n6503), .I1(n6122), .I2(n6507), .I3(n6123), 
            .O(n6508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__10199.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__10200 (.I0(\i16/rx_fifo/buff[23][3] ), .I1(\i16/rx_fifo/buff[21][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10200.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10201 (.I0(\i16/rx_fifo/buff[20][3] ), .I1(\i16/rx_fifo/buff[22][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10201.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10202 (.I0(\i16/rx_fifo/buff[19][3] ), .I1(\i16/rx_fifo/buff[17][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10202.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10203 (.I0(\i16/rx_fifo/buff[16][3] ), .I1(\i16/rx_fifo/buff[18][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10203.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10204 (.I0(n6512), .I1(n6122), .I2(n6511), .I3(n6123), 
            .O(n6513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10204.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10205 (.I0(n6509), .I1(n6510), .I2(n6122), .I3(n6513), 
            .O(n6514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10205.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10206 (.I0(n6508), .I1(n6514), .I2(n6127), .O(n6515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10206.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10207 (.I0(\i16/rx_fifo/buff[15][3] ), .I1(\i16/rx_fifo/buff[13][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10207.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10208 (.I0(\i16/rx_fifo/buff[12][3] ), .I1(\i16/rx_fifo/buff[14][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10208.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10209 (.I0(\i16/rx_fifo/buff[11][3] ), .I1(\i16/rx_fifo/buff[9][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10209.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10210 (.I0(\i16/rx_fifo/buff[8][3] ), .I1(\i16/rx_fifo/buff[10][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10210.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10211 (.I0(n6518), .I1(n6519), .I2(n6517), .I3(n6122), 
            .O(n6520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10211.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10212 (.I0(n6516), .I1(n6122), .I2(n6520), .I3(n6123), 
            .O(n6521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__10212.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__10213 (.I0(\i16/rx_fifo/buff[7][3] ), .I1(\i16/rx_fifo/buff[5][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10213.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10214 (.I0(\i16/rx_fifo/buff[4][3] ), .I1(\i16/rx_fifo/buff[6][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10214.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10215 (.I0(\i16/rx_fifo/buff[3][3] ), .I1(\i16/rx_fifo/buff[1][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10215.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10216 (.I0(\i16/rx_fifo/buff[0][3] ), .I1(\i16/rx_fifo/buff[2][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10216.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10217 (.I0(n6524), .I1(n6525), .I2(n6523), .I3(n6122), 
            .O(n6526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10217.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10218 (.I0(n6522), .I1(n6122), .I2(n6123), .I3(n6526), 
            .O(n6527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0c */ ;
    defparam LUT__10218.LUTMASK = 16'h0b0c;
    EFX_LUT4 LUT__10219 (.I0(n6521), .I1(n6127), .I2(n6527), .I3(n6117), 
            .O(n6528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10219.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10220 (.I0(\i16/rx_fifo/buff[39][3] ), .I1(\i16/rx_fifo/buff[37][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10220.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10221 (.I0(\i16/rx_fifo/buff[36][3] ), .I1(\i16/rx_fifo/buff[38][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10221.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10222 (.I0(\i16/rx_fifo/buff[35][3] ), .I1(\i16/rx_fifo/buff[33][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10222.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10223 (.I0(\i16/rx_fifo/buff[32][3] ), .I1(\i16/rx_fifo/buff[34][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10223.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10224 (.I0(n6531), .I1(n6532), .I2(n6530), .I3(n6122), 
            .O(n6533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10224.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10225 (.I0(n6529), .I1(n6122), .I2(n6123), .I3(n6533), 
            .O(n6534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0c */ ;
    defparam LUT__10225.LUTMASK = 16'h0b0c;
    EFX_LUT4 LUT__10226 (.I0(\i16/rx_fifo/buff[43][3] ), .I1(\i16/rx_fifo/buff[41][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10226.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10227 (.I0(\i16/rx_fifo/buff[40][3] ), .I1(\i16/rx_fifo/buff[42][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10227.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10228 (.I0(\i16/rx_fifo/buff[44][3] ), .I1(\i16/rx_fifo/buff[46][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10228.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10229 (.I0(n6535), .I1(n6536), .I2(n6537), .I3(n6122), 
            .O(n6538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10229.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10230 (.I0(\i16/rx_fifo/buff[47][3] ), .I1(\i16/rx_fifo/buff[45][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10230.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10231 (.I0(n6539), .I1(n6122), .I2(n6538), .I3(n6123), 
            .O(n6540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__10231.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__10232 (.I0(n6534), .I1(n6540), .I2(n6404), .O(n6541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10232.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10233 (.I0(\i16/rx_fifo/buff[51][3] ), .I1(\i16/rx_fifo/buff[49][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10233.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10234 (.I0(\i16/rx_fifo/buff[48][3] ), .I1(\i16/rx_fifo/buff[50][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10234.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10235 (.I0(n6542), .I1(n6543), .I2(n6122), .O(n6544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10235.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10236 (.I0(\i16/rx_fifo/buff[55][3] ), .I1(\i16/rx_fifo/buff[53][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10236.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10237 (.I0(\i16/rx_fifo/buff[52][3] ), .I1(\i16/rx_fifo/buff[54][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10237.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10238 (.I0(n6545), .I1(n6546), .I2(n6122), .I3(n6123), 
            .O(n6547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10238.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10239 (.I0(\i16/rx_fifo/buff[63][3] ), .I1(\i16/rx_fifo/buff[61][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10239.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10240 (.I0(\i16/rx_fifo/buff[60][3] ), .I1(\i16/rx_fifo/buff[62][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10240.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10241 (.I0(n6548), .I1(n6549), .I2(n6122), .O(n6550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10241.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10242 (.I0(\i16/rx_fifo/buff[59][3] ), .I1(\i16/rx_fifo/buff[57][3] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10242.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10243 (.I0(\i16/rx_fifo/buff[56][3] ), .I1(\i16/rx_fifo/buff[58][3] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10243.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10244 (.I0(n6552), .I1(n6122), .I2(n6551), .I3(n6123), 
            .O(n6553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10244.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10245 (.I0(n6550), .I1(n6553), .I2(n6544), .I3(n6547), 
            .O(n6554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10245.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10246 (.I0(n6405), .I1(n6554), .I2(n6119), .O(n6555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__10246.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__10247 (.I0(n6541), .I1(n6555), .I2(n6515), .I3(n6528), 
            .O(n6556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10247.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10248 (.I0(n6201), .I1(\rx_d[3] ), .I2(n6502), .I3(n6556), 
            .O(\rx_fifo/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__10248.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__10249 (.I0(\i16/rx_fifo/buff[75][4] ), .I1(\i16/rx_fifo/buff[73][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10249.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10250 (.I0(\i16/rx_fifo/buff[72][4] ), .I1(\i16/rx_fifo/buff[74][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10250.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10251 (.I0(n6557), .I1(n6558), .I2(n6122), .O(n6559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10251.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10252 (.I0(\i16/rx_fifo/buff[79][4] ), .I1(\i16/rx_fifo/buff[77][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10252.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10253 (.I0(\i16/rx_fifo/buff[76][4] ), .I1(\i16/rx_fifo/buff[78][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10253.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10254 (.I0(n6560), .I1(n6561), .I2(n6122), .I3(n6123), 
            .O(n6562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10254.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10255 (.I0(\i16/rx_fifo/buff[71][4] ), .I1(\i16/rx_fifo/buff[69][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10255.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10256 (.I0(\i16/rx_fifo/buff[68][4] ), .I1(\i16/rx_fifo/buff[70][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10256.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10257 (.I0(n6563), .I1(n6564), .I2(n6122), .O(n6565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10257.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10258 (.I0(\i16/rx_fifo/buff[67][4] ), .I1(\i16/rx_fifo/buff[65][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10258.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10259 (.I0(\i16/rx_fifo/buff[64][4] ), .I1(\i16/rx_fifo/buff[66][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10259.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10260 (.I0(n6567), .I1(n6122), .I2(n6566), .I3(n6123), 
            .O(n6568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10260.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10261 (.I0(n6565), .I1(n6568), .I2(n6559), .I3(n6562), 
            .O(n6569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10261.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10262 (.I0(\i16/rx_fifo/buff[111][4] ), .I1(\i16/rx_fifo/buff[109][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10262.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10263 (.I0(\i16/rx_fifo/buff[108][4] ), .I1(\i16/rx_fifo/buff[110][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10263.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10264 (.I0(n6570), .I1(n6571), .I2(n6122), .O(n6572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10264.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10265 (.I0(\i16/rx_fifo/buff[107][4] ), .I1(\i16/rx_fifo/buff[105][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10265.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10266 (.I0(\i16/rx_fifo/buff[104][4] ), .I1(\i16/rx_fifo/buff[106][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10266.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10267 (.I0(n6574), .I1(n6122), .I2(n6573), .I3(n6123), 
            .O(n6575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10267.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10268 (.I0(\i16/rx_fifo/buff[103][4] ), .I1(\i16/rx_fifo/buff[101][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10268.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10269 (.I0(\i16/rx_fifo/buff[100][4] ), .I1(\i16/rx_fifo/buff[102][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10269.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10270 (.I0(n6576), .I1(n6577), .I2(n6122), .O(n6578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10270.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10271 (.I0(\i16/rx_fifo/buff[99][4] ), .I1(\i16/rx_fifo/buff[97][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10271.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10272 (.I0(\i16/rx_fifo/buff[96][4] ), .I1(\i16/rx_fifo/buff[98][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10272.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10273 (.I0(n6580), .I1(n6122), .I2(n6579), .I3(n6123), 
            .O(n6581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10273.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10274 (.I0(n6578), .I1(n6581), .I2(n6572), .I3(n6575), 
            .O(n6582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10274.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10275 (.I0(n6582), .I1(n6569), .I2(n6127), .I3(n6117), 
            .O(n6583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10275.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10276 (.I0(\i16/rx_fifo/buff[119][4] ), .I1(\i16/rx_fifo/buff[117][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10276.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10277 (.I0(\i16/rx_fifo/buff[116][4] ), .I1(\i16/rx_fifo/buff[118][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10277.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10278 (.I0(n6584), .I1(n6585), .I2(n6122), .O(n6586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10278.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10279 (.I0(\i16/rx_fifo/buff[115][4] ), .I1(\i16/rx_fifo/buff[113][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10279.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10280 (.I0(\i16/rx_fifo/buff[112][4] ), .I1(\i16/rx_fifo/buff[114][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10280.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10281 (.I0(n6588), .I1(n6122), .I2(n6587), .I3(n6123), 
            .O(n6589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10281.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10282 (.I0(\i16/rx_fifo/buff[127][4] ), .I1(\i16/rx_fifo/buff[125][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10282.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10283 (.I0(\i16/rx_fifo/buff[124][4] ), .I1(\i16/rx_fifo/buff[126][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10283.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10284 (.I0(n6590), .I1(n6591), .I2(n6122), .O(n6592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10284.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10285 (.I0(\i16/rx_fifo/buff[123][4] ), .I1(\i16/rx_fifo/buff[121][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10285.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10286 (.I0(\i16/rx_fifo/buff[120][4] ), .I1(\i16/rx_fifo/buff[122][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10286.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10287 (.I0(n6594), .I1(n6122), .I2(n6593), .I3(n6123), 
            .O(n6595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10287.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10288 (.I0(n6592), .I1(n6595), .I2(n6586), .I3(n6589), 
            .O(n6596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10288.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10289 (.I0(\i16/rx_fifo/buff[83][4] ), .I1(\i16/rx_fifo/buff[81][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10289.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10290 (.I0(\i16/rx_fifo/buff[80][4] ), .I1(\i16/rx_fifo/buff[82][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10290.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10291 (.I0(n6597), .I1(n6598), .I2(n6122), .O(n6599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10291.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10292 (.I0(\i16/rx_fifo/buff[87][4] ), .I1(\i16/rx_fifo/buff[85][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10292.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10293 (.I0(\i16/rx_fifo/buff[84][4] ), .I1(\i16/rx_fifo/buff[86][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10293.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10294 (.I0(n6600), .I1(n6601), .I2(n6122), .I3(n6123), 
            .O(n6602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10294.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10295 (.I0(\i16/rx_fifo/buff[95][4] ), .I1(\i16/rx_fifo/buff[93][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10295.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10296 (.I0(\i16/rx_fifo/buff[92][4] ), .I1(\i16/rx_fifo/buff[94][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10296.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10297 (.I0(n6603), .I1(n6604), .I2(n6122), .O(n6605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10297.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10298 (.I0(\i16/rx_fifo/buff[91][4] ), .I1(\i16/rx_fifo/buff[89][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10298.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10299 (.I0(\i16/rx_fifo/buff[88][4] ), .I1(\i16/rx_fifo/buff[90][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10299.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10300 (.I0(n6607), .I1(n6122), .I2(n6606), .I3(n6123), 
            .O(n6608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10300.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10301 (.I0(n6605), .I1(n6608), .I2(n6599), .I3(n6602), 
            .O(n6609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10301.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10302 (.I0(n6609), .I1(n6596), .I2(\rx_fifo/rd_index[5] ), 
            .I3(n6127), .O(n6610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__10302.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__10303 (.I0(n6583), .I1(n6610), .I2(n6185), .O(n6611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10303.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10304 (.I0(\i16/rx_fifo/buff[31][4] ), .I1(\i16/rx_fifo/buff[29][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10304.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10305 (.I0(\i16/rx_fifo/buff[28][4] ), .I1(\i16/rx_fifo/buff[30][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10305.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10306 (.I0(\i16/rx_fifo/buff[27][4] ), .I1(\i16/rx_fifo/buff[25][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10306.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10307 (.I0(\i16/rx_fifo/buff[24][4] ), .I1(\i16/rx_fifo/buff[26][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10307.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10308 (.I0(n6614), .I1(n6615), .I2(n6613), .I3(n6122), 
            .O(n6616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10308.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10309 (.I0(n6612), .I1(n6122), .I2(n6616), .I3(n6123), 
            .O(n6617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__10309.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__10310 (.I0(\i16/rx_fifo/buff[23][4] ), .I1(\i16/rx_fifo/buff[21][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10310.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10311 (.I0(\i16/rx_fifo/buff[20][4] ), .I1(\i16/rx_fifo/buff[22][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6619)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10311.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10312 (.I0(\i16/rx_fifo/buff[19][4] ), .I1(\i16/rx_fifo/buff[17][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10312.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10313 (.I0(\i16/rx_fifo/buff[16][4] ), .I1(\i16/rx_fifo/buff[18][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6621)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10313.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10314 (.I0(n6621), .I1(n6122), .I2(n6620), .I3(n6123), 
            .O(n6622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10314.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10315 (.I0(n6618), .I1(n6619), .I2(n6122), .I3(n6622), 
            .O(n6623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10315.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10316 (.I0(n6617), .I1(n6623), .I2(n6127), .O(n6624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10316.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10317 (.I0(\i16/rx_fifo/buff[15][4] ), .I1(\i16/rx_fifo/buff[13][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10317.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10318 (.I0(\i16/rx_fifo/buff[12][4] ), .I1(\i16/rx_fifo/buff[14][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10318.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10319 (.I0(\i16/rx_fifo/buff[11][4] ), .I1(\i16/rx_fifo/buff[9][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10319.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10320 (.I0(\i16/rx_fifo/buff[8][4] ), .I1(\i16/rx_fifo/buff[10][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10320.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10321 (.I0(n6627), .I1(n6628), .I2(n6626), .I3(n6122), 
            .O(n6629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10321.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10322 (.I0(n6625), .I1(n6122), .I2(n6629), .I3(n6123), 
            .O(n6630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__10322.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__10323 (.I0(\i16/rx_fifo/buff[7][4] ), .I1(\i16/rx_fifo/buff[5][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10323.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10324 (.I0(\i16/rx_fifo/buff[4][4] ), .I1(\i16/rx_fifo/buff[6][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10324.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10325 (.I0(\i16/rx_fifo/buff[3][4] ), .I1(\i16/rx_fifo/buff[1][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10325.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10326 (.I0(\i16/rx_fifo/buff[0][4] ), .I1(\i16/rx_fifo/buff[2][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10326.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10327 (.I0(n6633), .I1(n6634), .I2(n6632), .I3(n6122), 
            .O(n6635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10327.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10328 (.I0(n6631), .I1(n6122), .I2(n6123), .I3(n6635), 
            .O(n6636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0c */ ;
    defparam LUT__10328.LUTMASK = 16'h0b0c;
    EFX_LUT4 LUT__10329 (.I0(n6630), .I1(n6127), .I2(n6636), .I3(n6117), 
            .O(n6637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10329.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10330 (.I0(\i16/rx_fifo/buff[39][4] ), .I1(\i16/rx_fifo/buff[37][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10330.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10331 (.I0(\i16/rx_fifo/buff[36][4] ), .I1(\i16/rx_fifo/buff[38][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10331.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10332 (.I0(\i16/rx_fifo/buff[35][4] ), .I1(\i16/rx_fifo/buff[33][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6640)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10332.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10333 (.I0(\i16/rx_fifo/buff[32][4] ), .I1(\i16/rx_fifo/buff[34][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10333.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10334 (.I0(n6640), .I1(n6641), .I2(n6639), .I3(n6122), 
            .O(n6642)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10334.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10335 (.I0(n6638), .I1(n6122), .I2(n6123), .I3(n6642), 
            .O(n6643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0c */ ;
    defparam LUT__10335.LUTMASK = 16'h0b0c;
    EFX_LUT4 LUT__10336 (.I0(\i16/rx_fifo/buff[43][4] ), .I1(\i16/rx_fifo/buff[41][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10336.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10337 (.I0(\i16/rx_fifo/buff[40][4] ), .I1(\i16/rx_fifo/buff[42][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10337.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10338 (.I0(\i16/rx_fifo/buff[44][4] ), .I1(\i16/rx_fifo/buff[46][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10338.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10339 (.I0(n6644), .I1(n6645), .I2(n6646), .I3(n6122), 
            .O(n6647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10339.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10340 (.I0(\i16/rx_fifo/buff[47][4] ), .I1(\i16/rx_fifo/buff[45][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10340.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10341 (.I0(n6648), .I1(n6122), .I2(n6647), .I3(n6123), 
            .O(n6649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__10341.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__10342 (.I0(n6643), .I1(n6649), .I2(n6404), .O(n6650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10342.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10343 (.I0(\i16/rx_fifo/buff[51][4] ), .I1(\i16/rx_fifo/buff[49][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10343.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10344 (.I0(\i16/rx_fifo/buff[48][4] ), .I1(\i16/rx_fifo/buff[50][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10344.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10345 (.I0(n6651), .I1(n6652), .I2(n6122), .O(n6653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10345.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10346 (.I0(\i16/rx_fifo/buff[55][4] ), .I1(\i16/rx_fifo/buff[53][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10346.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10347 (.I0(\i16/rx_fifo/buff[52][4] ), .I1(\i16/rx_fifo/buff[54][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10347.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10348 (.I0(n6654), .I1(n6655), .I2(n6122), .I3(n6123), 
            .O(n6656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10348.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10349 (.I0(\i16/rx_fifo/buff[63][4] ), .I1(\i16/rx_fifo/buff[61][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10349.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10350 (.I0(\i16/rx_fifo/buff[60][4] ), .I1(\i16/rx_fifo/buff[62][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10350.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10351 (.I0(n6657), .I1(n6658), .I2(n6122), .O(n6659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10351.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10352 (.I0(\i16/rx_fifo/buff[59][4] ), .I1(\i16/rx_fifo/buff[57][4] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10352.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10353 (.I0(\i16/rx_fifo/buff[56][4] ), .I1(\i16/rx_fifo/buff[58][4] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10353.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10354 (.I0(n6661), .I1(n6122), .I2(n6660), .I3(n6123), 
            .O(n6662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10354.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10355 (.I0(n6659), .I1(n6662), .I2(n6653), .I3(n6656), 
            .O(n6663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10355.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10356 (.I0(n6405), .I1(n6663), .I2(n6119), .O(n6664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__10356.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__10357 (.I0(n6650), .I1(n6664), .I2(n6624), .I3(n6637), 
            .O(n6665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10357.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10358 (.I0(n6201), .I1(\rx_d[4] ), .I2(n6611), .I3(n6665), 
            .O(\rx_fifo/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__10358.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__10359 (.I0(\i16/rx_fifo/buff[75][5] ), .I1(\i16/rx_fifo/buff[73][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10359.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10360 (.I0(\i16/rx_fifo/buff[72][5] ), .I1(\i16/rx_fifo/buff[74][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10360.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10361 (.I0(n6666), .I1(n6667), .I2(n6122), .O(n6668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10361.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10362 (.I0(\i16/rx_fifo/buff[79][5] ), .I1(\i16/rx_fifo/buff[77][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10362.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10363 (.I0(\i16/rx_fifo/buff[76][5] ), .I1(\i16/rx_fifo/buff[78][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10363.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10364 (.I0(n6669), .I1(n6670), .I2(n6122), .I3(n6123), 
            .O(n6671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10364.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10365 (.I0(\i16/rx_fifo/buff[71][5] ), .I1(\i16/rx_fifo/buff[69][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10365.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10366 (.I0(\i16/rx_fifo/buff[68][5] ), .I1(\i16/rx_fifo/buff[70][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10366.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10367 (.I0(n6672), .I1(n6673), .I2(n6122), .O(n6674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10367.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10368 (.I0(\i16/rx_fifo/buff[67][5] ), .I1(\i16/rx_fifo/buff[65][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10368.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10369 (.I0(\i16/rx_fifo/buff[64][5] ), .I1(\i16/rx_fifo/buff[66][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10369.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10370 (.I0(n6676), .I1(n6122), .I2(n6675), .I3(n6123), 
            .O(n6677)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10370.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10371 (.I0(n6674), .I1(n6677), .I2(n6668), .I3(n6671), 
            .O(n6678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10371.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10372 (.I0(\i16/rx_fifo/buff[111][5] ), .I1(\i16/rx_fifo/buff[109][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6679)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10372.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10373 (.I0(\i16/rx_fifo/buff[108][5] ), .I1(\i16/rx_fifo/buff[110][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10373.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10374 (.I0(n6679), .I1(n6680), .I2(n6122), .O(n6681)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10374.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10375 (.I0(\i16/rx_fifo/buff[107][5] ), .I1(\i16/rx_fifo/buff[105][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10375.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10376 (.I0(\i16/rx_fifo/buff[104][5] ), .I1(\i16/rx_fifo/buff[106][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10376.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10377 (.I0(n6683), .I1(n6122), .I2(n6682), .I3(n6123), 
            .O(n6684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10377.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10378 (.I0(\i16/rx_fifo/buff[103][5] ), .I1(\i16/rx_fifo/buff[101][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10378.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10379 (.I0(\i16/rx_fifo/buff[100][5] ), .I1(\i16/rx_fifo/buff[102][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10379.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10380 (.I0(n6685), .I1(n6686), .I2(n6122), .O(n6687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10380.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10381 (.I0(\i16/rx_fifo/buff[99][5] ), .I1(\i16/rx_fifo/buff[97][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10381.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10382 (.I0(\i16/rx_fifo/buff[96][5] ), .I1(\i16/rx_fifo/buff[98][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10382.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10383 (.I0(n6689), .I1(n6122), .I2(n6688), .I3(n6123), 
            .O(n6690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10383.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10384 (.I0(n6687), .I1(n6690), .I2(n6681), .I3(n6684), 
            .O(n6691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10384.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10385 (.I0(n6691), .I1(n6678), .I2(n6127), .I3(n6117), 
            .O(n6692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10385.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10386 (.I0(\i16/rx_fifo/buff[95][5] ), .I1(\i16/rx_fifo/buff[93][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10386.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10387 (.I0(\i16/rx_fifo/buff[92][5] ), .I1(\i16/rx_fifo/buff[94][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10387.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10388 (.I0(n6693), .I1(n6694), .I2(n6122), .O(n6695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10388.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10389 (.I0(\i16/rx_fifo/buff[91][5] ), .I1(\i16/rx_fifo/buff[89][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10389.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10390 (.I0(\i16/rx_fifo/buff[88][5] ), .I1(\i16/rx_fifo/buff[90][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10390.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10391 (.I0(n6697), .I1(n6122), .I2(n6696), .I3(n6123), 
            .O(n6698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10391.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10392 (.I0(\i16/rx_fifo/buff[83][5] ), .I1(\i16/rx_fifo/buff[81][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6699)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10392.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10393 (.I0(\i16/rx_fifo/buff[80][5] ), .I1(\i16/rx_fifo/buff[82][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6700)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10393.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10394 (.I0(n6699), .I1(n6700), .I2(n6122), .O(n6701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10394.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10395 (.I0(\i16/rx_fifo/buff[87][5] ), .I1(\i16/rx_fifo/buff[85][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6702)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10395.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10396 (.I0(\i16/rx_fifo/buff[84][5] ), .I1(\i16/rx_fifo/buff[86][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10396.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10397 (.I0(n6702), .I1(n6703), .I2(n6122), .I3(n6123), 
            .O(n6704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10397.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10398 (.I0(n6701), .I1(n6704), .I2(n6695), .I3(n6698), 
            .O(n6705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10398.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10399 (.I0(\i16/rx_fifo/buff[127][5] ), .I1(\i16/rx_fifo/buff[125][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10399.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10400 (.I0(\i16/rx_fifo/buff[124][5] ), .I1(\i16/rx_fifo/buff[126][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10400.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10401 (.I0(n6706), .I1(n6707), .I2(n6122), .O(n6708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10401.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10402 (.I0(\i16/rx_fifo/buff[123][5] ), .I1(\i16/rx_fifo/buff[121][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10402.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10403 (.I0(\i16/rx_fifo/buff[120][5] ), .I1(\i16/rx_fifo/buff[122][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10403.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10404 (.I0(n6710), .I1(n6122), .I2(n6709), .I3(n6123), 
            .O(n6711)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10404.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10405 (.I0(\i16/rx_fifo/buff[119][5] ), .I1(\i16/rx_fifo/buff[117][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6712)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10405.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10406 (.I0(\i16/rx_fifo/buff[116][5] ), .I1(\i16/rx_fifo/buff[118][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10406.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10407 (.I0(n6712), .I1(n6713), .I2(n6122), .O(n6714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10407.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10408 (.I0(\i16/rx_fifo/buff[115][5] ), .I1(\i16/rx_fifo/buff[113][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10408.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10409 (.I0(\i16/rx_fifo/buff[112][5] ), .I1(\i16/rx_fifo/buff[114][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10409.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10410 (.I0(n6716), .I1(n6122), .I2(n6715), .I3(n6123), 
            .O(n6717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10410.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10411 (.I0(n6714), .I1(n6717), .I2(n6708), .I3(n6711), 
            .O(n6718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10411.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10412 (.I0(n6718), .I1(n6705), .I2(\rx_fifo/rd_index[5] ), 
            .I3(n6127), .O(n6719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10412.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10413 (.I0(n6692), .I1(n6719), .I2(n6185), .O(n6720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10413.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10414 (.I0(\i16/rx_fifo/buff[55][5] ), .I1(\i16/rx_fifo/buff[53][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10414.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10415 (.I0(\i16/rx_fifo/buff[52][5] ), .I1(\i16/rx_fifo/buff[54][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10415.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10416 (.I0(\i16/rx_fifo/buff[48][5] ), .I1(\i16/rx_fifo/buff[50][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .O(n6723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10416.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10417 (.I0(\i16/rx_fifo/buff[51][5] ), .I1(\i16/rx_fifo/buff[49][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .O(n6724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__10417.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__10418 (.I0(n6724), .I1(n6723), .I2(n6122), .I3(\rx_fifo/rd_index[0] ), 
            .O(n6725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__10418.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__10419 (.I0(n6721), .I1(n6722), .I2(n6122), .I3(n6725), 
            .O(n6726)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10419.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10420 (.I0(\i16/rx_fifo/buff[59][5] ), .I1(\i16/rx_fifo/buff[57][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10420.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10421 (.I0(\i16/rx_fifo/buff[56][5] ), .I1(\i16/rx_fifo/buff[58][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10421.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10422 (.I0(\i16/rx_fifo/buff[60][5] ), .I1(\i16/rx_fifo/buff[62][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .O(n6729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10422.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10423 (.I0(\i16/rx_fifo/buff[63][5] ), .I1(\i16/rx_fifo/buff[61][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .O(n6730)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__10423.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__10424 (.I0(n6730), .I1(n6729), .I2(\rx_fifo/rd_index[0] ), 
            .I3(n6122), .O(n6731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__10424.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__10425 (.I0(n6728), .I1(n6122), .I2(n6727), .I3(n6731), 
            .O(n6732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10425.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10426 (.I0(n6732), .I1(n6726), .I2(n6123), .O(n6733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10426.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10427 (.I0(\i16/rx_fifo/buff[43][5] ), .I1(\i16/rx_fifo/buff[41][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10427.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10428 (.I0(\i16/rx_fifo/buff[40][5] ), .I1(\i16/rx_fifo/buff[42][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10428.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10429 (.I0(\i16/rx_fifo/buff[47][5] ), .I1(\i16/rx_fifo/buff[45][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10429.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10430 (.I0(\i16/rx_fifo/buff[44][5] ), .I1(\i16/rx_fifo/buff[46][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10430.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10431 (.I0(n6736), .I1(n6737), .I2(n6122), .I3(n6123), 
            .O(n6738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10431.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10432 (.I0(n6735), .I1(n6122), .I2(n6734), .I3(n6738), 
            .O(n6739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10432.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10433 (.I0(\i16/rx_fifo/buff[39][5] ), .I1(\i16/rx_fifo/buff[37][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10433.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10434 (.I0(\i16/rx_fifo/buff[36][5] ), .I1(\i16/rx_fifo/buff[38][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10434.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10435 (.I0(\i16/rx_fifo/buff[35][5] ), .I1(\i16/rx_fifo/buff[33][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10435.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10436 (.I0(\i16/rx_fifo/buff[32][5] ), .I1(\i16/rx_fifo/buff[34][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10436.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10437 (.I0(n6743), .I1(n6122), .I2(n6742), .I3(n6123), 
            .O(n6744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10437.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10438 (.I0(n6740), .I1(n6741), .I2(n6122), .I3(n6744), 
            .O(n6745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10438.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10439 (.I0(n6745), .I1(n6739), .I2(n6404), .I3(n6119), 
            .O(n6746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10439.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10440 (.I0(\i16/rx_fifo/buff[7][5] ), .I1(\i16/rx_fifo/buff[5][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10440.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10441 (.I0(\i16/rx_fifo/buff[4][5] ), .I1(\i16/rx_fifo/buff[6][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10441.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10442 (.I0(n6747), .I1(n6748), .I2(n6122), .O(n6749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10442.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10443 (.I0(\i16/rx_fifo/buff[3][5] ), .I1(\i16/rx_fifo/buff[1][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10443.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10444 (.I0(\i16/rx_fifo/buff[0][5] ), .I1(\i16/rx_fifo/buff[2][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10444.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10445 (.I0(n6751), .I1(n6122), .I2(n6750), .I3(n6123), 
            .O(n6752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10445.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10446 (.I0(\i16/rx_fifo/buff[15][5] ), .I1(\i16/rx_fifo/buff[13][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10446.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10447 (.I0(\i16/rx_fifo/buff[12][5] ), .I1(\i16/rx_fifo/buff[14][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10447.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10448 (.I0(n6753), .I1(n6754), .I2(n6122), .O(n6755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10448.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10449 (.I0(\i16/rx_fifo/buff[11][5] ), .I1(\i16/rx_fifo/buff[9][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10449.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10450 (.I0(\i16/rx_fifo/buff[8][5] ), .I1(\i16/rx_fifo/buff[10][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10450.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10451 (.I0(n6757), .I1(n6122), .I2(n6756), .I3(n6123), 
            .O(n6758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10451.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10452 (.I0(n6755), .I1(n6758), .I2(n6749), .I3(n6752), 
            .O(n6759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10452.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10453 (.I0(\i16/rx_fifo/buff[31][5] ), .I1(\i16/rx_fifo/buff[29][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10453.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10454 (.I0(\i16/rx_fifo/buff[28][5] ), .I1(\i16/rx_fifo/buff[30][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10454.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10455 (.I0(n6760), .I1(n6761), .I2(n6122), .O(n6762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10455.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10456 (.I0(\i16/rx_fifo/buff[27][5] ), .I1(\i16/rx_fifo/buff[25][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10456.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10457 (.I0(\i16/rx_fifo/buff[24][5] ), .I1(\i16/rx_fifo/buff[26][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10457.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10458 (.I0(n6764), .I1(n6122), .I2(n6763), .I3(n6123), 
            .O(n6765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10458.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10459 (.I0(\i16/rx_fifo/buff[23][5] ), .I1(\i16/rx_fifo/buff[21][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6766)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10459.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10460 (.I0(\i16/rx_fifo/buff[20][5] ), .I1(\i16/rx_fifo/buff[22][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10460.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10461 (.I0(n6766), .I1(n6767), .I2(n6122), .O(n6768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10461.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10462 (.I0(\i16/rx_fifo/buff[19][5] ), .I1(\i16/rx_fifo/buff[17][5] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10462.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10463 (.I0(\i16/rx_fifo/buff[16][5] ), .I1(\i16/rx_fifo/buff[18][5] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10463.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10464 (.I0(n6770), .I1(n6122), .I2(n6769), .I3(n6123), 
            .O(n6771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10464.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10465 (.I0(n6768), .I1(n6771), .I2(n6762), .I3(n6765), 
            .O(n6772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10465.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10466 (.I0(n6772), .I1(n6759), .I2(n6117), .I3(n6127), 
            .O(n6773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10466.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10467 (.I0(n6405), .I1(n6733), .I2(n6746), .I3(n6773), 
            .O(n6774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__10467.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__10468 (.I0(n6201), .I1(\rx_d[5] ), .I2(n6720), .I3(n6774), 
            .O(\rx_fifo/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__10468.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__10469 (.I0(\i16/rx_fifo/buff[116][6] ), .I1(\i16/rx_fifo/buff[118][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10469.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10470 (.I0(\i16/rx_fifo/buff[117][6] ), .I1(\i16/rx_fifo/buff[119][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6775), .O(n6776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc */ ;
    defparam LUT__10470.LUTMASK = 16'h0afc;
    EFX_LUT4 LUT__10471 (.I0(\i16/rx_fifo/buff[112][6] ), .I1(\i16/rx_fifo/buff[114][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10471.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10472 (.I0(\i16/rx_fifo/buff[115][6] ), .I1(\i16/rx_fifo/buff[113][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6777), .O(n6778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10472.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10473 (.I0(n6778), .I1(n6776), .I2(n6123), .I3(n6122), 
            .O(n6779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__10473.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__10474 (.I0(\i16/rx_fifo/buff[123][6] ), .I1(\i16/rx_fifo/buff[121][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10474.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10475 (.I0(\i16/rx_fifo/buff[120][6] ), .I1(\i16/rx_fifo/buff[122][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10475.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10476 (.I0(\i16/rx_fifo/buff[127][6] ), .I1(\i16/rx_fifo/buff[125][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10476.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10477 (.I0(\i16/rx_fifo/buff[124][6] ), .I1(\i16/rx_fifo/buff[126][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10477.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10478 (.I0(n6782), .I1(n6783), .I2(n6122), .I3(n6123), 
            .O(n6784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10478.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10479 (.I0(n6781), .I1(n6122), .I2(n6780), .I3(n6784), 
            .O(n6785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10479.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10480 (.I0(\i16/rx_fifo/buff[87][6] ), .I1(\i16/rx_fifo/buff[85][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10480.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10481 (.I0(\i16/rx_fifo/buff[84][6] ), .I1(\i16/rx_fifo/buff[86][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10481.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10482 (.I0(n6786), .I1(n6787), .I2(n6122), .O(n6788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10482.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10483 (.I0(\i16/rx_fifo/buff[83][6] ), .I1(\i16/rx_fifo/buff[81][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10483.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10484 (.I0(\i16/rx_fifo/buff[80][6] ), .I1(\i16/rx_fifo/buff[82][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10484.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10485 (.I0(n6790), .I1(n6122), .I2(n6789), .I3(n6123), 
            .O(n6791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10485.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10486 (.I0(\i16/rx_fifo/buff[91][6] ), .I1(\i16/rx_fifo/buff[89][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10486.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10487 (.I0(\i16/rx_fifo/buff[88][6] ), .I1(\i16/rx_fifo/buff[90][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10487.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10488 (.I0(n6792), .I1(n6793), .I2(n6122), .O(n6794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10488.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10489 (.I0(\i16/rx_fifo/buff[95][6] ), .I1(\i16/rx_fifo/buff[93][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10489.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10490 (.I0(\i16/rx_fifo/buff[92][6] ), .I1(\i16/rx_fifo/buff[94][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10490.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10491 (.I0(n6795), .I1(n6796), .I2(n6122), .I3(n6123), 
            .O(n6797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10491.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10492 (.I0(n6794), .I1(n6797), .I2(n6788), .I3(n6791), 
            .O(n6798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10492.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10493 (.I0(n6785), .I1(n6779), .I2(n6798), .I3(n6117), 
            .O(n6799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__10493.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__10494 (.I0(n6799), .I1(n6127), .I2(n6185), .O(n6800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__10494.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__10495 (.I0(\i16/rx_fifo/buff[103][6] ), .I1(\i16/rx_fifo/buff[101][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10495.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10496 (.I0(\rx_fifo/rd_index[1] ), .I1(\i16/rx_fifo/buff[102][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .O(n6802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10496.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10497 (.I0(\rx_fifo/rd_index[2] ), .I1(\i16/rx_fifo/buff[100][6] ), 
            .I2(n6801), .I3(n6802), .O(n6803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__10497.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__10498 (.I0(\i16/rx_fifo/buff[96][6] ), .I1(\i16/rx_fifo/buff[98][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10498.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10499 (.I0(\i16/rx_fifo/buff[99][6] ), .I1(\i16/rx_fifo/buff[97][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6804), .O(n6805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10499.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10500 (.I0(n6803), .I1(n6805), .I2(n6123), .I3(n6122), 
            .O(n6806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05fc */ ;
    defparam LUT__10500.LUTMASK = 16'h05fc;
    EFX_LUT4 LUT__10501 (.I0(\i16/rx_fifo/buff[111][6] ), .I1(\i16/rx_fifo/buff[109][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10501.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10502 (.I0(\i16/rx_fifo/buff[108][6] ), .I1(\i16/rx_fifo/buff[110][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10502.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10503 (.I0(\i16/rx_fifo/buff[107][6] ), .I1(\i16/rx_fifo/buff[105][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10503.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10504 (.I0(\i16/rx_fifo/buff[104][6] ), .I1(\i16/rx_fifo/buff[106][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10504.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10505 (.I0(n6809), .I1(n6810), .I2(n6808), .I3(n6122), 
            .O(n6811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__10505.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__10506 (.I0(n6807), .I1(n6806), .I2(n6811), .I3(n6123), 
            .O(n6812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d33 */ ;
    defparam LUT__10506.LUTMASK = 16'h0d33;
    EFX_LUT4 LUT__10507 (.I0(\i16/rx_fifo/buff[75][6] ), .I1(\i16/rx_fifo/buff[73][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10507.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10508 (.I0(\i16/rx_fifo/buff[72][6] ), .I1(\i16/rx_fifo/buff[74][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6814)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10508.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10509 (.I0(\i16/rx_fifo/buff[76][6] ), .I1(\i16/rx_fifo/buff[78][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10509.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10510 (.I0(n6813), .I1(n6814), .I2(n6815), .I3(n6122), 
            .O(n6816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__10510.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__10511 (.I0(\i16/rx_fifo/buff[79][6] ), .I1(\i16/rx_fifo/buff[77][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10511.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10512 (.I0(\i16/rx_fifo/buff[71][6] ), .I1(\i16/rx_fifo/buff[69][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10512.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10513 (.I0(\i16/rx_fifo/buff[68][6] ), .I1(\i16/rx_fifo/buff[70][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10513.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10514 (.I0(n6818), .I1(n6819), .I2(n6817), .I3(n6123), 
            .O(n6820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10514.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10515 (.I0(\i16/rx_fifo/buff[67][6] ), .I1(\i16/rx_fifo/buff[65][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10515.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10516 (.I0(\i16/rx_fifo/buff[64][6] ), .I1(\i16/rx_fifo/buff[66][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10516.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10517 (.I0(n6821), .I1(n6822), .I2(n6820), .I3(n6122), 
            .O(n6823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__10517.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__10518 (.I0(n6122), .I1(n6816), .I2(n6123), .I3(n6823), 
            .O(n6824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h301f */ ;
    defparam LUT__10518.LUTMASK = 16'h301f;
    EFX_LUT4 LUT__10519 (.I0(n6824), .I1(n6812), .I2(n6127), .I3(n6117), 
            .O(n6825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__10519.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__10520 (.I0(\i16/rx_fifo/buff[39][6] ), .I1(\i16/rx_fifo/buff[37][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10520.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10521 (.I0(\i16/rx_fifo/buff[36][6] ), .I1(\i16/rx_fifo/buff[38][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10521.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10522 (.I0(\i16/rx_fifo/buff[32][6] ), .I1(\i16/rx_fifo/buff[34][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10522.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10523 (.I0(\i16/rx_fifo/buff[35][6] ), .I1(\i16/rx_fifo/buff[33][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6828), .O(n6829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10523.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10524 (.I0(n6827), .I1(n6826), .I2(n6829), .I3(n6122), 
            .O(n6830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10524.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10525 (.I0(\i16/rx_fifo/buff[47][6] ), .I1(\i16/rx_fifo/buff[45][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10525.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10526 (.I0(\i16/rx_fifo/buff[44][6] ), .I1(\i16/rx_fifo/buff[46][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10526.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10527 (.I0(\i16/rx_fifo/buff[43][6] ), .I1(\i16/rx_fifo/buff[41][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10527.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10528 (.I0(\i16/rx_fifo/buff[40][6] ), .I1(\i16/rx_fifo/buff[42][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10528.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10529 (.I0(n6833), .I1(n6834), .I2(n6122), .O(n6835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10529.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10530 (.I0(n6831), .I1(n6832), .I2(n6122), .I3(n6835), 
            .O(n6836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10530.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10531 (.I0(n6836), .I1(n6830), .I2(n6127), .I3(n6123), 
            .O(n6837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10531.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10532 (.I0(\i16/rx_fifo/buff[63][6] ), .I1(\i16/rx_fifo/buff[61][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10532.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10533 (.I0(\i16/rx_fifo/buff[60][6] ), .I1(\i16/rx_fifo/buff[62][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10533.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10534 (.I0(\i16/rx_fifo/buff[59][6] ), .I1(\i16/rx_fifo/buff[57][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10534.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10535 (.I0(\i16/rx_fifo/buff[56][6] ), .I1(\i16/rx_fifo/buff[58][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10535.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10536 (.I0(n6840), .I1(n6841), .I2(n6839), .I3(n6122), 
            .O(n6842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10536.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10537 (.I0(n6838), .I1(n6122), .I2(n6842), .I3(n6123), 
            .O(n6843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__10537.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__10538 (.I0(\i16/rx_fifo/buff[48][6] ), .I1(\i16/rx_fifo/buff[50][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10538.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10539 (.I0(\i16/rx_fifo/buff[51][6] ), .I1(\i16/rx_fifo/buff[49][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6844), .O(n6845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10539.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10540 (.I0(\i16/rx_fifo/buff[55][6] ), .I1(\i16/rx_fifo/buff[53][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10540.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10541 (.I0(\rx_fifo/rd_index[1] ), .I1(\i16/rx_fifo/buff[54][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .O(n6847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10541.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10542 (.I0(\rx_fifo/rd_index[2] ), .I1(\i16/rx_fifo/buff[52][6] ), 
            .I2(n6846), .I3(n6847), .O(n6848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__10542.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__10543 (.I0(n6848), .I1(n6845), .I2(n6123), .I3(n6122), 
            .O(n6849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__10543.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__10544 (.I0(n6843), .I1(n6849), .I2(n6127), .I3(n6117), 
            .O(n6850)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10544.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10545 (.I0(\i16/rx_fifo/buff[7][6] ), .I1(\i16/rx_fifo/buff[5][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10545.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10546 (.I0(\i16/rx_fifo/buff[4][6] ), .I1(\i16/rx_fifo/buff[6][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10546.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10547 (.I0(\i16/rx_fifo/buff[3][6] ), .I1(\i16/rx_fifo/buff[1][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10547.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10548 (.I0(\i16/rx_fifo/buff[0][6] ), .I1(\i16/rx_fifo/buff[2][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10548.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10549 (.I0(n6853), .I1(n6854), .I2(n6122), .O(n6855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10549.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10550 (.I0(n6851), .I1(n6852), .I2(n6122), .I3(n6855), 
            .O(n6856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10550.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10551 (.I0(\i16/rx_fifo/buff[15][6] ), .I1(\i16/rx_fifo/buff[13][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10551.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10552 (.I0(\i16/rx_fifo/buff[12][6] ), .I1(\i16/rx_fifo/buff[14][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10552.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10553 (.I0(\i16/rx_fifo/buff[11][6] ), .I1(\i16/rx_fifo/buff[9][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10553.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10554 (.I0(\i16/rx_fifo/buff[8][6] ), .I1(\i16/rx_fifo/buff[10][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10554.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10555 (.I0(n6859), .I1(n6860), .I2(n6122), .O(n6861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10555.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10556 (.I0(n6857), .I1(n6858), .I2(n6122), .I3(n6861), 
            .O(n6862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10556.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10557 (.I0(n6862), .I1(n6856), .I2(n6123), .I3(n6404), 
            .O(n6863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10557.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10558 (.I0(\i16/rx_fifo/buff[23][6] ), .I1(\i16/rx_fifo/buff[21][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10558.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10559 (.I0(\i16/rx_fifo/buff[20][6] ), .I1(\i16/rx_fifo/buff[22][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10559.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10560 (.I0(\i16/rx_fifo/buff[19][6] ), .I1(\i16/rx_fifo/buff[17][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10560.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10561 (.I0(\i16/rx_fifo/buff[16][6] ), .I1(\i16/rx_fifo/buff[18][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10561.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10562 (.I0(n6866), .I1(n6867), .I2(n6865), .I3(n6122), 
            .O(n6868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10562.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10563 (.I0(n6864), .I1(n6122), .I2(n6123), .I3(n6868), 
            .O(n6869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0c */ ;
    defparam LUT__10563.LUTMASK = 16'h0b0c;
    EFX_LUT4 LUT__10564 (.I0(\i16/rx_fifo/buff[31][6] ), .I1(\i16/rx_fifo/buff[29][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10564.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10565 (.I0(\i16/rx_fifo/buff[28][6] ), .I1(\i16/rx_fifo/buff[30][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10565.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10566 (.I0(\i16/rx_fifo/buff[27][6] ), .I1(\i16/rx_fifo/buff[25][6] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10566.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10567 (.I0(\i16/rx_fifo/buff[24][6] ), .I1(\i16/rx_fifo/buff[26][6] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10567.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10568 (.I0(n6873), .I1(n6122), .I2(n6872), .I3(n6123), 
            .O(n6874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10568.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10569 (.I0(n6870), .I1(n6871), .I2(n6122), .I3(n6874), 
            .O(n6875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10569.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10570 (.I0(n6875), .I1(n6869), .I2(n6405), .I3(n6227), 
            .O(n6876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10570.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10571 (.I0(n6863), .I1(n6876), .I2(n6837), .I3(n6850), 
            .O(n6877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10571.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10572 (.I0(n6201), .I1(\rx_d[6] ), .O(n6878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10572.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10573 (.I0(n6825), .I1(n6800), .I2(n6877), .I3(n6878), 
            .O(\rx_fifo/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4 */ ;
    defparam LUT__10573.LUTMASK = 16'hfff4;
    EFX_LUT4 LUT__10574 (.I0(\i16/rx_fifo/buff[71][7] ), .I1(\i16/rx_fifo/buff[69][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10574.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10575 (.I0(\i16/rx_fifo/buff[68][7] ), .I1(\i16/rx_fifo/buff[70][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10575.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10576 (.I0(\i16/rx_fifo/buff[67][7] ), .I1(\i16/rx_fifo/buff[65][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10576.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10577 (.I0(\i16/rx_fifo/buff[64][7] ), .I1(\i16/rx_fifo/buff[66][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10577.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10578 (.I0(n6881), .I1(n6882), .I2(n6122), .O(n6883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10578.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10579 (.I0(n6879), .I1(n6880), .I2(n6122), .I3(n6883), 
            .O(n6884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10579.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10580 (.I0(\i16/rx_fifo/buff[79][7] ), .I1(\i16/rx_fifo/buff[77][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10580.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10581 (.I0(\i16/rx_fifo/buff[76][7] ), .I1(\i16/rx_fifo/buff[78][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10581.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10582 (.I0(\i16/rx_fifo/buff[75][7] ), .I1(\i16/rx_fifo/buff[73][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10582.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10583 (.I0(\i16/rx_fifo/buff[72][7] ), .I1(\i16/rx_fifo/buff[74][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10583.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10584 (.I0(n6887), .I1(n6888), .I2(n6122), .O(n6889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10584.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10585 (.I0(n6885), .I1(n6886), .I2(n6122), .I3(n6889), 
            .O(n6890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10585.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10586 (.I0(n6890), .I1(n6884), .I2(n6117), .I3(n6123), 
            .O(n6891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10586.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10587 (.I0(\i16/rx_fifo/buff[103][7] ), .I1(\i16/rx_fifo/buff[101][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10587.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10588 (.I0(\i16/rx_fifo/buff[100][7] ), .I1(\i16/rx_fifo/buff[102][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10588.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10589 (.I0(\i16/rx_fifo/buff[99][7] ), .I1(\i16/rx_fifo/buff[97][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10589.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10590 (.I0(\i16/rx_fifo/buff[96][7] ), .I1(\i16/rx_fifo/buff[98][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10590.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10591 (.I0(n6894), .I1(n6895), .I2(n6122), .O(n6896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10591.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10592 (.I0(n6892), .I1(n6893), .I2(n6122), .I3(n6896), 
            .O(n6897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10592.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10593 (.I0(\i16/rx_fifo/buff[111][7] ), .I1(\i16/rx_fifo/buff[109][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10593.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10594 (.I0(\i16/rx_fifo/buff[108][7] ), .I1(\i16/rx_fifo/buff[110][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10594.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10595 (.I0(\i16/rx_fifo/buff[104][7] ), .I1(\i16/rx_fifo/buff[106][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10595.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10596 (.I0(\i16/rx_fifo/buff[107][7] ), .I1(\i16/rx_fifo/buff[105][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6900), .O(n6901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10596.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10597 (.I0(n6899), .I1(n6898), .I2(n6901), .I3(n6122), 
            .O(n6902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10597.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10598 (.I0(n6902), .I1(n6897), .I2(n6123), .I3(n6117), 
            .O(n6903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10598.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10599 (.I0(\i16/rx_fifo/buff[112][7] ), .I1(\i16/rx_fifo/buff[114][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10599.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10600 (.I0(\i16/rx_fifo/buff[115][7] ), .I1(\i16/rx_fifo/buff[113][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6904), .O(n6905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10600.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10601 (.I0(\i16/rx_fifo/buff[119][7] ), .I1(\i16/rx_fifo/buff[117][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10601.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10602 (.I0(\rx_fifo/rd_index[1] ), .I1(\i16/rx_fifo/buff[118][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .O(n6907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10602.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10603 (.I0(\rx_fifo/rd_index[2] ), .I1(\i16/rx_fifo/buff[116][7] ), 
            .I2(n6906), .I3(n6907), .O(n6908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__10603.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__10604 (.I0(n6908), .I1(n6905), .I2(n6123), .I3(n6122), 
            .O(n6909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__10604.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__10605 (.I0(\i16/rx_fifo/buff[120][7] ), .I1(\i16/rx_fifo/buff[122][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10605.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10606 (.I0(\i16/rx_fifo/buff[123][7] ), .I1(\i16/rx_fifo/buff[121][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6910), .O(n6911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10606.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10607 (.I0(\i16/rx_fifo/buff[127][7] ), .I1(\i16/rx_fifo/buff[125][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10607.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10608 (.I0(\i16/rx_fifo/buff[124][7] ), .I1(\i16/rx_fifo/buff[126][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10608.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10609 (.I0(n6912), .I1(n6913), .I2(n6122), .I3(n6123), 
            .O(n6914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10609.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10610 (.I0(n6122), .I1(n6911), .I2(n6914), .I3(n6117), 
            .O(n6915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__10610.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__10611 (.I0(\i16/rx_fifo/buff[87][7] ), .I1(\i16/rx_fifo/buff[85][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10611.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10612 (.I0(\rx_fifo/rd_index[1] ), .I1(\i16/rx_fifo/buff[86][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .O(n6917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10612.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10613 (.I0(\rx_fifo/rd_index[2] ), .I1(\i16/rx_fifo/buff[84][7] ), 
            .I2(n6916), .I3(n6917), .O(n6918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__10613.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__10614 (.I0(\i16/rx_fifo/buff[80][7] ), .I1(\i16/rx_fifo/buff[82][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10614.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10615 (.I0(\i16/rx_fifo/buff[83][7] ), .I1(\i16/rx_fifo/buff[81][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6919), .O(n6920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10615.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10616 (.I0(n6920), .I1(n6918), .I2(n6123), .I3(n6122), 
            .O(n6921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a */ ;
    defparam LUT__10616.LUTMASK = 16'h030a;
    EFX_LUT4 LUT__10617 (.I0(\i16/rx_fifo/buff[92][7] ), .I1(\i16/rx_fifo/buff[94][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10617.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10618 (.I0(\i16/rx_fifo/buff[95][7] ), .I1(\i16/rx_fifo/buff[93][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6922), .O(n6923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10618.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10619 (.I0(\i16/rx_fifo/buff[91][7] ), .I1(\i16/rx_fifo/buff[89][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10619.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10620 (.I0(\i16/rx_fifo/buff[88][7] ), .I1(\i16/rx_fifo/buff[90][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10620.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10621 (.I0(n6925), .I1(n6122), .I2(n6924), .I3(n6123), 
            .O(n6926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10621.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10622 (.I0(n6923), .I1(n6122), .I2(n6926), .I3(n6117), 
            .O(n6927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__10622.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__10623 (.I0(n6921), .I1(n6927), .I2(n6909), .I3(n6915), 
            .O(n6928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10623.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10624 (.I0(n6903), .I1(n6891), .I2(n6928), .I3(n6127), 
            .O(n6929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10624.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10625 (.I0(n6201), .I1(\rx_d[7] ), .O(n6930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10625.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10626 (.I0(\i16/rx_fifo/buff[39][7] ), .I1(\i16/rx_fifo/buff[37][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10626.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10627 (.I0(\i16/rx_fifo/buff[36][7] ), .I1(\i16/rx_fifo/buff[38][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10627.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10628 (.I0(\i16/rx_fifo/buff[35][7] ), .I1(\i16/rx_fifo/buff[33][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10628.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10629 (.I0(\i16/rx_fifo/buff[32][7] ), .I1(\i16/rx_fifo/buff[34][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10629.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10630 (.I0(n6934), .I1(n6122), .I2(n6933), .I3(n6123), 
            .O(n6935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10630.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10631 (.I0(n6931), .I1(n6932), .I2(n6122), .I3(n6935), 
            .O(n6936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10631.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10632 (.I0(\i16/rx_fifo/buff[47][7] ), .I1(\i16/rx_fifo/buff[45][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10632.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10633 (.I0(\i16/rx_fifo/buff[44][7] ), .I1(\i16/rx_fifo/buff[46][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10633.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10634 (.I0(\i16/rx_fifo/buff[43][7] ), .I1(\i16/rx_fifo/buff[41][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10634.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10635 (.I0(\i16/rx_fifo/buff[40][7] ), .I1(\i16/rx_fifo/buff[42][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10635.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10636 (.I0(n6940), .I1(n6122), .I2(n6939), .I3(n6123), 
            .O(n6941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10636.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10637 (.I0(n6937), .I1(n6938), .I2(n6122), .I3(n6941), 
            .O(n6942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10637.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10638 (.I0(n6936), .I1(n6942), .I2(n6127), .O(n6943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10638.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10639 (.I0(\i16/rx_fifo/buff[51][7] ), .I1(\i16/rx_fifo/buff[49][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10639.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10640 (.I0(\i16/rx_fifo/buff[48][7] ), .I1(\i16/rx_fifo/buff[50][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10640.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10641 (.I0(\i16/rx_fifo/buff[55][7] ), .I1(\i16/rx_fifo/buff[53][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10641.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10642 (.I0(\i16/rx_fifo/buff[52][7] ), .I1(\i16/rx_fifo/buff[54][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10642.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10643 (.I0(n6946), .I1(n6947), .I2(n6122), .I3(n6123), 
            .O(n6948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10643.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10644 (.I0(n6945), .I1(n6122), .I2(n6944), .I3(n6948), 
            .O(n6949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10644.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10645 (.I0(\i16/rx_fifo/buff[63][7] ), .I1(\i16/rx_fifo/buff[61][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10645.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10646 (.I0(\i16/rx_fifo/buff[60][7] ), .I1(\i16/rx_fifo/buff[62][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10646.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10647 (.I0(\i16/rx_fifo/buff[59][7] ), .I1(\i16/rx_fifo/buff[57][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10647.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10648 (.I0(\i16/rx_fifo/buff[56][7] ), .I1(\i16/rx_fifo/buff[58][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10648.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10649 (.I0(n6953), .I1(n6122), .I2(n6952), .I3(n6123), 
            .O(n6954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10649.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10650 (.I0(n6950), .I1(n6951), .I2(n6122), .I3(n6954), 
            .O(n6955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10650.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10651 (.I0(n6955), .I1(n6949), .I2(n6127), .I3(n6117), 
            .O(n6956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10651.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10652 (.I0(\i16/rx_fifo/buff[7][7] ), .I1(\i16/rx_fifo/buff[5][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10652.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10653 (.I0(\i16/rx_fifo/buff[4][7] ), .I1(\i16/rx_fifo/buff[6][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10653.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10654 (.I0(\i16/rx_fifo/buff[0][7] ), .I1(\i16/rx_fifo/buff[2][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10654.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10655 (.I0(\i16/rx_fifo/buff[3][7] ), .I1(\i16/rx_fifo/buff[1][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(n6959), .O(n6960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10655.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10656 (.I0(n6958), .I1(n6957), .I2(n6960), .I3(n6122), 
            .O(n6961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10656.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10657 (.I0(\i16/rx_fifo/buff[11][7] ), .I1(\i16/rx_fifo/buff[9][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10657.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10658 (.I0(\i16/rx_fifo/buff[8][7] ), .I1(\i16/rx_fifo/buff[10][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10658.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10659 (.I0(\i16/rx_fifo/buff[15][7] ), .I1(\i16/rx_fifo/buff[13][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10659.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10660 (.I0(\i16/rx_fifo/buff[12][7] ), .I1(\i16/rx_fifo/buff[14][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10660.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10661 (.I0(n6964), .I1(n6965), .I2(n6122), .I3(n6123), 
            .O(n6966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10661.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10662 (.I0(n6963), .I1(n6122), .I2(n6962), .I3(n6966), 
            .O(n6967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10662.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10663 (.I0(n6961), .I1(n6123), .I2(n6967), .I3(n6404), 
            .O(n6968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__10663.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__10664 (.I0(\i16/rx_fifo/buff[23][7] ), .I1(\i16/rx_fifo/buff[21][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10664.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10665 (.I0(\i16/rx_fifo/buff[20][7] ), .I1(\i16/rx_fifo/buff[22][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10665.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10666 (.I0(\i16/rx_fifo/buff[19][7] ), .I1(\i16/rx_fifo/buff[17][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10666.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10667 (.I0(\i16/rx_fifo/buff[16][7] ), .I1(\i16/rx_fifo/buff[18][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10667.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10668 (.I0(n6972), .I1(n6122), .I2(n6971), .I3(n6123), 
            .O(n6973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10668.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10669 (.I0(n6969), .I1(n6970), .I2(n6122), .I3(n6973), 
            .O(n6974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10669.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10670 (.I0(\i16/rx_fifo/buff[31][7] ), .I1(\i16/rx_fifo/buff[29][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10670.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10671 (.I0(\i16/rx_fifo/buff[28][7] ), .I1(\i16/rx_fifo/buff[30][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10671.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10672 (.I0(\i16/rx_fifo/buff[27][7] ), .I1(\i16/rx_fifo/buff[25][7] ), 
            .I2(\rx_fifo/rd_index[0] ), .I3(\rx_fifo/rd_index[1] ), .O(n6977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10672.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10673 (.I0(\i16/rx_fifo/buff[24][7] ), .I1(\i16/rx_fifo/buff[26][7] ), 
            .I2(\rx_fifo/rd_index[1] ), .I3(\rx_fifo/rd_index[0] ), .O(n6978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10673.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10674 (.I0(n6978), .I1(n6122), .I2(n6977), .I3(n6123), 
            .O(n6979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10674.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10675 (.I0(n6975), .I1(n6976), .I2(n6122), .I3(n6979), 
            .O(n6980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10675.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10676 (.I0(n6980), .I1(n6974), .I2(n6405), .I3(n6227), 
            .O(n6981)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10676.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10677 (.I0(n6968), .I1(n6981), .I2(n6943), .I3(n6956), 
            .O(n6982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__10677.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__10678 (.I0(n6929), .I1(n6185), .I2(n6930), .I3(n6982), 
            .O(\rx_fifo/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__10678.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__10679 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[3] ), 
            .I2(\fifo_inst/wr_index[4] ), .I3(\fifo_inst/wr_index[2] ), 
            .O(n6983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10679.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10680 (.I0(n4324), .I1(n6983), .O(\i14/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10680.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10681 (.I0(n4321), .I1(n6983), .O(\i14/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10681.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10682 (.I0(\fifo_inst/wr_index[3] ), .I1(\fifo_inst/wr_index[4] ), 
            .I2(\fifo_inst/wr_index[1] ), .I3(\fifo_inst/wr_index[2] ), 
            .O(n6984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10682.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10683 (.I0(n4324), .I1(n6984), .O(\i14/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10683.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10684 (.I0(n4321), .I1(n6984), .O(\i14/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10684.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10685 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[2] ), 
            .I2(\fifo_inst/wr_index[4] ), .I3(\fifo_inst/wr_index[3] ), 
            .O(n6985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10685.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10686 (.I0(n4324), .I1(n6985), .O(\i14/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10686.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10687 (.I0(n4321), .I1(n6985), .O(\i14/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10687.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10688 (.I0(\fifo_inst/wr_index[2] ), .I1(\fifo_inst/wr_index[4] ), 
            .I2(\fifo_inst/wr_index[3] ), .I3(\fifo_inst/wr_index[1] ), 
            .O(n6986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10688.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10689 (.I0(n4324), .I1(n6986), .O(\i14/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10689.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10690 (.I0(n4321), .I1(n6986), .O(\i14/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10690.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10691 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[4] ), 
            .I2(\fifo_inst/wr_index[3] ), .I3(\fifo_inst/wr_index[2] ), 
            .O(n6987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10691.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10692 (.I0(n4324), .I1(n6987), .O(\i14/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10692.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10693 (.I0(n4321), .I1(n6987), .O(\i14/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10693.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10694 (.I0(\fifo_inst/wr_index[4] ), .I1(\fifo_inst/wr_index[2] ), 
            .I2(\fifo_inst/wr_index[3] ), .I3(\fifo_inst/wr_index[1] ), 
            .O(n6988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10694.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10695 (.I0(n4324), .I1(n6988), .O(\i14/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10695.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10696 (.I0(n4321), .I1(n6988), .O(\i14/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10696.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10697 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[2] ), 
            .I2(\fifo_inst/wr_index[3] ), .I3(\fifo_inst/wr_index[4] ), 
            .O(n6989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10697.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10698 (.I0(n4324), .I1(n6989), .O(\i14/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10698.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10699 (.I0(n4321), .I1(n6989), .O(\i14/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10699.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10700 (.I0(\fifo_inst/wr_index[2] ), .I1(\fifo_inst/wr_index[3] ), 
            .I2(\fifo_inst/wr_index[1] ), .I3(\fifo_inst/wr_index[4] ), 
            .O(n6990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10700.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10701 (.I0(n4324), .I1(n6990), .O(\i14/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10701.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10702 (.I0(n4321), .I1(n6990), .O(\i14/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10702.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10703 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[3] ), 
            .I2(\fifo_inst/wr_index[2] ), .I3(\fifo_inst/wr_index[4] ), 
            .O(n6991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10703.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10704 (.I0(n4324), .I1(n6991), .O(\i14/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10704.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10705 (.I0(n4321), .I1(n6991), .O(\i14/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10705.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10706 (.I0(\fifo_inst/wr_index[3] ), .I1(\fifo_inst/wr_index[2] ), 
            .I2(\fifo_inst/wr_index[1] ), .I3(\fifo_inst/wr_index[4] ), 
            .O(n6992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10706.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10707 (.I0(n4324), .I1(n6992), .O(\i14/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10707.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10708 (.I0(n4321), .I1(n6992), .O(\i14/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10708.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10709 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[2] ), 
            .I2(\fifo_inst/wr_index[3] ), .I3(\fifo_inst/wr_index[4] ), 
            .O(n6993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10709.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10710 (.I0(n4324), .I1(n6993), .O(\i14/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10710.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10711 (.I0(n4321), .I1(n6993), .O(\i14/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10711.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10712 (.I0(\fifo_inst/wr_index[2] ), .I1(\fifo_inst/wr_index[1] ), 
            .I2(\fifo_inst/wr_index[3] ), .I3(\fifo_inst/wr_index[4] ), 
            .O(n6994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10712.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10713 (.I0(n4324), .I1(n6994), .O(\i14/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10713.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10714 (.I0(n4321), .I1(n6994), .O(\i14/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10714.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10715 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[2] ), 
            .I2(\fifo_inst/wr_index[3] ), .I3(\fifo_inst/wr_index[4] ), 
            .O(n6995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10715.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10716 (.I0(n4324), .I1(n6995), .O(\i14/n104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10716.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10717 (.I0(n4321), .I1(n6995), .O(\i14/n103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10717.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10718 (.I0(\fifo_inst/wr_index[1] ), .I1(\fifo_inst/wr_index[2] ), 
            .I2(\fifo_inst/wr_index[3] ), .I3(\fifo_inst/wr_index[4] ), 
            .O(n6996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10718.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10719 (.I0(n4324), .I1(n6996), .O(\i14/n102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10719.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10720 (.I0(n4321), .I1(n6996), .O(\i14/n101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10720.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10721 (.I0(\fifo_inst/wr_index[6] ), .I1(\fifo_inst/wr_index[5] ), 
            .I2(n4323), .O(n6997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10721.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10722 (.I0(n6997), .I1(n4476), .O(\i14/n100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10722.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10723 (.I0(\fifo_inst/wr_index[6] ), .I1(\fifo_inst/wr_index[5] ), 
            .I2(n4320), .O(n6998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10723.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10724 (.I0(n6998), .I1(n4476), .O(\i14/n99 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10724.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10725 (.I0(n6997), .I1(n4322), .O(\i14/n98 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10725.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10726 (.I0(n6998), .I1(n4322), .O(\i14/n97 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10726.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10727 (.I0(n6997), .I1(n6983), .O(\i14/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10727.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10728 (.I0(n6998), .I1(n6983), .O(\i14/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10728.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10729 (.I0(n6997), .I1(n6984), .O(\i14/n94 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10729.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10730 (.I0(n6998), .I1(n6984), .O(\i14/n93 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10730.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10731 (.I0(n6997), .I1(n6985), .O(\i14/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10731.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10732 (.I0(n6998), .I1(n6985), .O(\i14/n91 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10732.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10733 (.I0(n6997), .I1(n6986), .O(\i14/n90 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10733.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10734 (.I0(n6998), .I1(n6986), .O(\i14/n89 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10734.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10735 (.I0(n6997), .I1(n6987), .O(\i14/n88 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10735.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10736 (.I0(n6998), .I1(n6987), .O(\i14/n87 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10736.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10737 (.I0(n6997), .I1(n6988), .O(\i14/n86 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10737.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10738 (.I0(n6998), .I1(n6988), .O(\i14/n85 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10738.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10739 (.I0(n6997), .I1(n6989), .O(\i14/n84 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10739.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10740 (.I0(n6998), .I1(n6989), .O(\i14/n83 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10740.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10741 (.I0(n6997), .I1(n6990), .O(\i14/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10741.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10742 (.I0(n6998), .I1(n6990), .O(\i14/n81 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10742.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10743 (.I0(n6997), .I1(n6991), .O(\i14/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10743.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10744 (.I0(n6998), .I1(n6991), .O(\i14/n79 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10744.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10745 (.I0(n6997), .I1(n6992), .O(\i14/n78 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10745.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10746 (.I0(n6998), .I1(n6992), .O(\i14/n77 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10746.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10747 (.I0(n6997), .I1(n6993), .O(\i14/n76 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10747.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10748 (.I0(n6998), .I1(n6993), .O(\i14/n75 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10748.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10749 (.I0(n6997), .I1(n6994), .O(\i14/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10749.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10750 (.I0(n6998), .I1(n6994), .O(\i14/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10750.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10751 (.I0(n6997), .I1(n6995), .O(\i14/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10751.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10752 (.I0(n6998), .I1(n6995), .O(\i14/n71 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10752.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10753 (.I0(n6997), .I1(n6996), .O(\i14/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10753.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10754 (.I0(n6998), .I1(n6996), .O(\i14/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10754.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10755 (.I0(\fifo_inst/wr_index[5] ), .I1(n4323), .I2(\fifo_inst/wr_index[6] ), 
            .O(n6999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10755.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10756 (.I0(n6999), .I1(n4476), .O(\i14/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10756.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10757 (.I0(\fifo_inst/wr_index[5] ), .I1(n4320), .I2(\fifo_inst/wr_index[6] ), 
            .O(n7000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10757.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10758 (.I0(n7000), .I1(n4476), .O(\i14/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10758.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10759 (.I0(n6999), .I1(n4322), .O(\i14/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10759.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10760 (.I0(n7000), .I1(n4322), .O(\i14/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10760.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10761 (.I0(n6999), .I1(n6983), .O(\i14/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10761.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10762 (.I0(n7000), .I1(n6983), .O(\i14/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10762.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10763 (.I0(n6999), .I1(n6984), .O(\i14/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10763.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10764 (.I0(n7000), .I1(n6984), .O(\i14/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10764.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10765 (.I0(n6999), .I1(n6985), .O(\i14/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10765.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10766 (.I0(n7000), .I1(n6985), .O(\i14/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10766.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10767 (.I0(n6999), .I1(n6986), .O(\i14/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10767.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10768 (.I0(n7000), .I1(n6986), .O(\i14/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10768.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10769 (.I0(n6999), .I1(n6987), .O(\i14/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10769.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10770 (.I0(n7000), .I1(n6987), .O(\i14/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10770.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10771 (.I0(n6999), .I1(n6988), .O(\i14/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10771.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10772 (.I0(n7000), .I1(n6988), .O(\i14/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10772.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10773 (.I0(n6999), .I1(n6989), .O(\i14/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10773.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10774 (.I0(n7000), .I1(n6989), .O(\i14/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10774.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10775 (.I0(n6999), .I1(n6990), .O(\i14/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10775.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10776 (.I0(n7000), .I1(n6990), .O(\i14/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10776.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10777 (.I0(n6999), .I1(n6991), .O(\i14/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10777.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10778 (.I0(n7000), .I1(n6991), .O(\i14/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10778.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10779 (.I0(n6999), .I1(n6992), .O(\i14/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10779.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10780 (.I0(n7000), .I1(n6992), .O(\i14/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10780.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10781 (.I0(n6999), .I1(n6993), .O(\i14/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10781.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10782 (.I0(n7000), .I1(n6993), .O(\i14/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10782.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10783 (.I0(n6999), .I1(n6994), .O(\i14/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10783.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10784 (.I0(n7000), .I1(n6994), .O(\i14/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10784.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10785 (.I0(n6999), .I1(n6995), .O(\i14/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10785.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10786 (.I0(n7000), .I1(n6995), .O(\i14/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10786.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10787 (.I0(n6999), .I1(n6996), .O(\i14/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10787.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10788 (.I0(n7000), .I1(n6996), .O(\i14/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10788.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10789 (.I0(n4323), .I1(\fifo_inst/wr_index[5] ), .I2(\fifo_inst/wr_index[6] ), 
            .O(n7001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10789.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10790 (.I0(n7001), .I1(n4476), .O(\i14/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10790.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10791 (.I0(n4320), .I1(\fifo_inst/wr_index[5] ), .I2(\fifo_inst/wr_index[6] ), 
            .O(n7002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10791.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10792 (.I0(n7002), .I1(n4476), .O(\i14/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10792.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10793 (.I0(n7001), .I1(n4322), .O(\i14/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10793.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10794 (.I0(n7002), .I1(n4322), .O(\i14/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10794.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10795 (.I0(n7001), .I1(n6983), .O(\i14/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10795.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10796 (.I0(n7002), .I1(n6983), .O(\i14/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10796.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10797 (.I0(n7001), .I1(n6984), .O(\i14/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10797.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10798 (.I0(n7002), .I1(n6984), .O(\i14/n29 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10798.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10799 (.I0(n7001), .I1(n6985), .O(\i14/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10799.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10800 (.I0(n7002), .I1(n6985), .O(\i14/n27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10800.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10801 (.I0(n7001), .I1(n6986), .O(\i14/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10801.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10802 (.I0(n7002), .I1(n6986), .O(\i14/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10802.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10803 (.I0(n7001), .I1(n6987), .O(\i14/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10803.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10804 (.I0(n7002), .I1(n6987), .O(\i14/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10804.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10805 (.I0(n7001), .I1(n6988), .O(\i14/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10805.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10806 (.I0(n7002), .I1(n6988), .O(\i14/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10806.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10807 (.I0(n7001), .I1(n6989), .O(\i14/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10807.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10808 (.I0(n7002), .I1(n6989), .O(\i14/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10808.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10809 (.I0(n7001), .I1(n6990), .O(\i14/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10809.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10810 (.I0(n7002), .I1(n6990), .O(\i14/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10810.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10811 (.I0(n7001), .I1(n6991), .O(\i14/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10811.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10812 (.I0(n7002), .I1(n6991), .O(\i14/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10812.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10813 (.I0(n7001), .I1(n6992), .O(\i14/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10813.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10814 (.I0(n7002), .I1(n6992), .O(\i14/n13 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10814.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10815 (.I0(n7001), .I1(n6993), .O(\i14/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10815.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10816 (.I0(n7002), .I1(n6993), .O(\i14/n11 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10816.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10817 (.I0(n7001), .I1(n6994), .O(\i14/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10817.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10818 (.I0(n7002), .I1(n6994), .O(\i14/n9 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10818.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10819 (.I0(n7001), .I1(n6995), .O(\i14/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10819.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10820 (.I0(n7002), .I1(n6995), .O(\i14/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10820.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10821 (.I0(n7001), .I1(n6996), .O(\i14/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10821.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10822 (.I0(n7002), .I1(n6996), .O(\i14/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10822.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10823 (.I0(\tx_fifo/wr_index[0] ), .I1(\tx_fifo/wr_index[7] ), 
            .I2(n5232), .O(n7003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10823.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10824 (.I0(\tx_fifo/wr_index[5] ), .I1(\tx_fifo/wr_index[6] ), 
            .I2(n7003), .O(n7004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10824.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10825 (.I0(\tx_fifo/wr_index[1] ), .I1(\tx_fifo/wr_index[2] ), 
            .I2(\tx_fifo/wr_index[3] ), .I3(\tx_fifo/wr_index[4] ), .O(n7005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10825.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10826 (.I0(n7004), .I1(n7005), .O(\i15/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10826.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10827 (.I0(\tx_fifo/wr_index[7] ), .I1(\tx_fifo/wr_index[0] ), 
            .I2(n5232), .O(n7006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10827.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10828 (.I0(\tx_fifo/wr_index[5] ), .I1(\tx_fifo/wr_index[6] ), 
            .I2(n7006), .O(n7007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10828.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10829 (.I0(n7007), .I1(n7005), .O(\i15/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10829.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10830 (.I0(\tx_fifo/wr_index[2] ), .I1(\tx_fifo/wr_index[3] ), 
            .I2(\tx_fifo/wr_index[4] ), .I3(\tx_fifo/wr_index[1] ), .O(n7008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10830.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10831 (.I0(n7004), .I1(n7008), .O(\i15/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10831.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10832 (.I0(n7007), .I1(n7008), .O(\i15/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10832.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10833 (.I0(\tx_fifo/wr_index[1] ), .I1(\tx_fifo/wr_index[3] ), 
            .I2(\tx_fifo/wr_index[4] ), .I3(\tx_fifo/wr_index[2] ), .O(n7009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10833.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10834 (.I0(n7004), .I1(n7009), .O(\i15/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10834.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10835 (.I0(n7007), .I1(n7009), .O(\i15/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10835.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10836 (.I0(\tx_fifo/wr_index[3] ), .I1(\tx_fifo/wr_index[4] ), 
            .I2(\tx_fifo/wr_index[1] ), .I3(\tx_fifo/wr_index[2] ), .O(n7010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10836.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10837 (.I0(n7004), .I1(n7010), .O(\i15/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10837.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10838 (.I0(n7007), .I1(n7010), .O(\i15/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10838.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10839 (.I0(\tx_fifo/wr_index[1] ), .I1(\tx_fifo/wr_index[2] ), 
            .I2(\tx_fifo/wr_index[4] ), .I3(\tx_fifo/wr_index[3] ), .O(n7011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10839.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10840 (.I0(n7004), .I1(n7011), .O(\i15/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10840.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10841 (.I0(n7007), .I1(n7011), .O(\i15/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10841.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10842 (.I0(\tx_fifo/wr_index[2] ), .I1(\tx_fifo/wr_index[4] ), 
            .I2(\tx_fifo/wr_index[3] ), .I3(\tx_fifo/wr_index[1] ), .O(n7012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10842.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10843 (.I0(n7004), .I1(n7012), .O(\i15/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10843.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10844 (.I0(n7007), .I1(n7012), .O(\i15/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10844.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10845 (.I0(\tx_fifo/wr_index[1] ), .I1(\tx_fifo/wr_index[4] ), 
            .I2(\tx_fifo/wr_index[3] ), .I3(\tx_fifo/wr_index[2] ), .O(n7013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10845.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10846 (.I0(n7004), .I1(n7013), .O(\i15/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10846.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10847 (.I0(n7007), .I1(n7013), .O(\i15/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10847.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10848 (.I0(\tx_fifo/wr_index[4] ), .I1(\tx_fifo/wr_index[2] ), 
            .I2(\tx_fifo/wr_index[3] ), .I3(\tx_fifo/wr_index[1] ), .O(n7014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10848.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10849 (.I0(n7004), .I1(n7014), .O(\i15/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10849.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10850 (.I0(n7007), .I1(n7014), .O(\i15/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10850.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10851 (.I0(\tx_fifo/wr_index[1] ), .I1(\tx_fifo/wr_index[2] ), 
            .I2(\tx_fifo/wr_index[3] ), .I3(\tx_fifo/wr_index[4] ), .O(n7015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10851.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10852 (.I0(n7004), .I1(n7015), .O(\i15/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10852.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10853 (.I0(n7007), .I1(n7015), .O(\i15/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10853.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10854 (.I0(\tx_fifo/wr_index[2] ), .I1(\tx_fifo/wr_index[3] ), 
            .I2(\tx_fifo/wr_index[1] ), .I3(\tx_fifo/wr_index[4] ), .O(n7016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10854.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10855 (.I0(n7004), .I1(n7016), .O(\i15/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10855.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10856 (.I0(n7007), .I1(n7016), .O(\i15/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10856.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10857 (.I0(\tx_fifo/wr_index[1] ), .I1(\tx_fifo/wr_index[3] ), 
            .I2(\tx_fifo/wr_index[2] ), .I3(\tx_fifo/wr_index[4] ), .O(n7017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10857.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10858 (.I0(n7004), .I1(n7017), .O(\i15/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10858.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10859 (.I0(n7007), .I1(n7017), .O(\i15/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10859.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10860 (.I0(\tx_fifo/wr_index[3] ), .I1(\tx_fifo/wr_index[2] ), 
            .I2(\tx_fifo/wr_index[1] ), .I3(\tx_fifo/wr_index[4] ), .O(n7018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10860.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10861 (.I0(n7004), .I1(n7018), .O(\i15/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10861.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10862 (.I0(n7007), .I1(n7018), .O(\i15/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10862.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10863 (.I0(\tx_fifo/wr_index[1] ), .I1(\tx_fifo/wr_index[2] ), 
            .I2(\tx_fifo/wr_index[3] ), .I3(\tx_fifo/wr_index[4] ), .O(n7019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10863.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10864 (.I0(n7004), .I1(n7019), .O(\i15/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10864.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10865 (.I0(n7007), .I1(n7019), .O(\i15/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10865.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10866 (.I0(\tx_fifo/wr_index[2] ), .I1(\tx_fifo/wr_index[1] ), 
            .I2(\tx_fifo/wr_index[3] ), .I3(\tx_fifo/wr_index[4] ), .O(n7020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10866.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10867 (.I0(n7004), .I1(n7020), .O(\i15/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10867.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10868 (.I0(n7007), .I1(n7020), .O(\i15/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10868.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10869 (.I0(\tx_fifo/wr_index[1] ), .I1(\tx_fifo/wr_index[2] ), 
            .I2(\tx_fifo/wr_index[3] ), .I3(\tx_fifo/wr_index[4] ), .O(n7021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10869.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10870 (.I0(n7004), .I1(n7021), .O(\i15/n104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10870.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10871 (.I0(n7007), .I1(n7021), .O(\i15/n103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10871.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10872 (.I0(\tx_fifo/wr_index[1] ), .I1(\tx_fifo/wr_index[2] ), 
            .I2(\tx_fifo/wr_index[3] ), .I3(\tx_fifo/wr_index[4] ), .O(n7022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10872.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10873 (.I0(n7004), .I1(n7022), .O(\i15/n102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10873.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10874 (.I0(n7007), .I1(n7022), .O(\i15/n101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10874.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10875 (.I0(\tx_fifo/wr_index[6] ), .I1(\tx_fifo/wr_index[5] ), 
            .I2(n7003), .O(n7023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10875.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10876 (.I0(n7023), .I1(n7005), .O(\i15/n100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10876.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10877 (.I0(\tx_fifo/wr_index[6] ), .I1(\tx_fifo/wr_index[5] ), 
            .I2(n7006), .O(n7024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10877.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10878 (.I0(n7024), .I1(n7005), .O(\i15/n99 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10878.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10879 (.I0(n7023), .I1(n7008), .O(\i15/n98 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10879.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10880 (.I0(n7024), .I1(n7008), .O(\i15/n97 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10880.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10881 (.I0(n7023), .I1(n7009), .O(\i15/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10881.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10882 (.I0(n7024), .I1(n7009), .O(\i15/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10882.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10883 (.I0(n7023), .I1(n7010), .O(\i15/n94 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10883.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10884 (.I0(n7024), .I1(n7010), .O(\i15/n93 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10884.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10885 (.I0(n7023), .I1(n7011), .O(\i15/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10885.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10886 (.I0(n7024), .I1(n7011), .O(\i15/n91 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10886.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10887 (.I0(n7023), .I1(n7012), .O(\i15/n90 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10887.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10888 (.I0(n7024), .I1(n7012), .O(\i15/n89 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10888.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10889 (.I0(n7023), .I1(n7013), .O(\i15/n88 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10889.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10890 (.I0(n7024), .I1(n7013), .O(\i15/n87 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10890.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10891 (.I0(n7023), .I1(n7014), .O(\i15/n86 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10891.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10892 (.I0(n7024), .I1(n7014), .O(\i15/n85 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10892.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10893 (.I0(n7023), .I1(n7015), .O(\i15/n84 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10893.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10894 (.I0(n7024), .I1(n7015), .O(\i15/n83 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10894.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10895 (.I0(n7023), .I1(n7016), .O(\i15/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10895.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10896 (.I0(n7024), .I1(n7016), .O(\i15/n81 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10896.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10897 (.I0(n7023), .I1(n7017), .O(\i15/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10897.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10898 (.I0(n7024), .I1(n7017), .O(\i15/n79 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10898.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10899 (.I0(n7023), .I1(n7018), .O(\i15/n78 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10899.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10900 (.I0(n7024), .I1(n7018), .O(\i15/n77 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10900.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10901 (.I0(n7023), .I1(n7019), .O(\i15/n76 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10901.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10902 (.I0(n7024), .I1(n7019), .O(\i15/n75 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10902.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10903 (.I0(n7023), .I1(n7020), .O(\i15/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10903.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10904 (.I0(n7024), .I1(n7020), .O(\i15/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10904.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10905 (.I0(n7023), .I1(n7021), .O(\i15/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10905.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10906 (.I0(n7024), .I1(n7021), .O(\i15/n71 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10906.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10907 (.I0(n7023), .I1(n7022), .O(\i15/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10907.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10908 (.I0(n7024), .I1(n7022), .O(\i15/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10908.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10909 (.I0(\tx_fifo/wr_index[5] ), .I1(n7003), .I2(\tx_fifo/wr_index[6] ), 
            .O(n7025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10909.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10910 (.I0(n7025), .I1(n7005), .O(\i15/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10910.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10911 (.I0(\tx_fifo/wr_index[5] ), .I1(n7006), .I2(\tx_fifo/wr_index[6] ), 
            .O(n7026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10911.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10912 (.I0(n7026), .I1(n7005), .O(\i15/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10912.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10913 (.I0(n7025), .I1(n7008), .O(\i15/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10913.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10914 (.I0(n7026), .I1(n7008), .O(\i15/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10914.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10915 (.I0(n7025), .I1(n7009), .O(\i15/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10915.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10916 (.I0(n7026), .I1(n7009), .O(\i15/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10916.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10917 (.I0(n7025), .I1(n7010), .O(\i15/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10917.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10918 (.I0(n7026), .I1(n7010), .O(\i15/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10918.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10919 (.I0(n7025), .I1(n7011), .O(\i15/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10919.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10920 (.I0(n7026), .I1(n7011), .O(\i15/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10920.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10921 (.I0(n7025), .I1(n7012), .O(\i15/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10921.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10922 (.I0(n7026), .I1(n7012), .O(\i15/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10922.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10923 (.I0(n7025), .I1(n7013), .O(\i15/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10923.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10924 (.I0(n7026), .I1(n7013), .O(\i15/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10924.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10925 (.I0(n7025), .I1(n7014), .O(\i15/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10925.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10926 (.I0(n7026), .I1(n7014), .O(\i15/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10926.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10927 (.I0(n7025), .I1(n7015), .O(\i15/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10927.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10928 (.I0(n7026), .I1(n7015), .O(\i15/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10928.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10929 (.I0(n7025), .I1(n7016), .O(\i15/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10929.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10930 (.I0(n7026), .I1(n7016), .O(\i15/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10930.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10931 (.I0(n7025), .I1(n7017), .O(\i15/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10931.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10932 (.I0(n7026), .I1(n7017), .O(\i15/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10932.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10933 (.I0(n7025), .I1(n7018), .O(\i15/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10933.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10934 (.I0(n7026), .I1(n7018), .O(\i15/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10934.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10935 (.I0(n7025), .I1(n7019), .O(\i15/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10935.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10936 (.I0(n7026), .I1(n7019), .O(\i15/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10936.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10937 (.I0(n7025), .I1(n7020), .O(\i15/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10937.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10938 (.I0(n7026), .I1(n7020), .O(\i15/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10938.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10939 (.I0(n7025), .I1(n7021), .O(\i15/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10939.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10940 (.I0(n7026), .I1(n7021), .O(\i15/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10940.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10941 (.I0(n7025), .I1(n7022), .O(\i15/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10941.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10942 (.I0(n7026), .I1(n7022), .O(\i15/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10942.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10943 (.I0(n7003), .I1(\tx_fifo/wr_index[5] ), .I2(\tx_fifo/wr_index[6] ), 
            .O(n7027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10943.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10944 (.I0(n7027), .I1(n7005), .O(\i15/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10944.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10945 (.I0(n7006), .I1(\tx_fifo/wr_index[5] ), .I2(\tx_fifo/wr_index[6] ), 
            .O(n7028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10945.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10946 (.I0(n7028), .I1(n7005), .O(\i15/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10946.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10947 (.I0(n7027), .I1(n7008), .O(\i15/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10947.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10948 (.I0(n7028), .I1(n7008), .O(\i15/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10948.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10949 (.I0(n7027), .I1(n7009), .O(\i15/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10949.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10950 (.I0(n7028), .I1(n7009), .O(\i15/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10950.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10951 (.I0(n7027), .I1(n7010), .O(\i15/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10951.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10952 (.I0(n7028), .I1(n7010), .O(\i15/n29 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10952.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10953 (.I0(n7027), .I1(n7011), .O(\i15/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10953.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10954 (.I0(n7028), .I1(n7011), .O(\i15/n27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10954.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10955 (.I0(n7027), .I1(n7012), .O(\i15/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10955.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10956 (.I0(n7028), .I1(n7012), .O(\i15/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10956.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10957 (.I0(n7027), .I1(n7013), .O(\i15/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10957.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10958 (.I0(n7028), .I1(n7013), .O(\i15/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10958.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10959 (.I0(n7027), .I1(n7014), .O(\i15/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10959.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10960 (.I0(n7028), .I1(n7014), .O(\i15/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10960.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10961 (.I0(n7027), .I1(n7015), .O(\i15/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10961.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10962 (.I0(n7028), .I1(n7015), .O(\i15/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10962.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10963 (.I0(n7027), .I1(n7016), .O(\i15/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10963.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10964 (.I0(n7028), .I1(n7016), .O(\i15/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10964.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10965 (.I0(n7027), .I1(n7017), .O(\i15/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10965.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10966 (.I0(n7028), .I1(n7017), .O(\i15/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10966.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10967 (.I0(n7027), .I1(n7018), .O(\i15/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10967.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10968 (.I0(n7028), .I1(n7018), .O(\i15/n13 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10968.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10969 (.I0(n7027), .I1(n7019), .O(\i15/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10969.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10970 (.I0(n7028), .I1(n7019), .O(\i15/n11 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10970.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10971 (.I0(n7027), .I1(n7020), .O(\i15/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10971.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10972 (.I0(n7028), .I1(n7020), .O(\i15/n9 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10972.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10973 (.I0(n7027), .I1(n7021), .O(\i15/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10973.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10974 (.I0(n7028), .I1(n7021), .O(\i15/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10974.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10975 (.I0(n7027), .I1(n7022), .O(\i15/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10975.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10976 (.I0(n7028), .I1(n7022), .O(\i15/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10976.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10977 (.I0(rx_en_rx_packet), .I1(\rx_d[0] ), .O(\data_to_rx_packet_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10977.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10978 (.I0(\rx_fifo/wr_index[0] ), .I1(\rx_fifo/wr_index[7] ), 
            .I2(n6109), .O(n7029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10978.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10979 (.I0(\rx_fifo/wr_index[5] ), .I1(\rx_fifo/wr_index[6] ), 
            .I2(n7029), .O(n7030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10979.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10980 (.I0(\rx_fifo/wr_index[1] ), .I1(\rx_fifo/wr_index[2] ), 
            .I2(\rx_fifo/wr_index[3] ), .I3(\rx_fifo/wr_index[4] ), .O(n7031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10980.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10981 (.I0(n7030), .I1(n7031), .O(\i16/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10981.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10982 (.I0(rx_en_rx_packet), .I1(\rx_d[1] ), .O(\data_to_rx_packet_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10982.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10983 (.I0(rx_en_rx_packet), .I1(\rx_d[2] ), .O(\data_to_rx_packet_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10983.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10984 (.I0(rx_en_rx_packet), .I1(\rx_d[3] ), .O(\data_to_rx_packet_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10984.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10985 (.I0(rx_en_rx_packet), .I1(\rx_d[4] ), .O(\data_to_rx_packet_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10985.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10986 (.I0(rx_en_rx_packet), .I1(\rx_d[5] ), .O(\data_to_rx_packet_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10986.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10987 (.I0(rx_en_rx_packet), .I1(\rx_d[6] ), .O(\data_to_rx_packet_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10987.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10988 (.I0(rx_en_rx_packet), .I1(\rx_d[7] ), .O(\data_to_rx_packet_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10988.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10989 (.I0(\rx_fifo/wr_index[7] ), .I1(\rx_fifo/wr_index[0] ), 
            .I2(n6109), .O(n7032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10989.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10990 (.I0(\rx_fifo/wr_index[5] ), .I1(\rx_fifo/wr_index[6] ), 
            .I2(n7032), .O(n7033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10990.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10991 (.I0(n7033), .I1(n7031), .O(\i16/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10991.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10992 (.I0(\rx_fifo/wr_index[2] ), .I1(\rx_fifo/wr_index[3] ), 
            .I2(\rx_fifo/wr_index[4] ), .I3(\rx_fifo/wr_index[1] ), .O(n7034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10992.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10993 (.I0(n7030), .I1(n7034), .O(\i16/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10993.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10994 (.I0(n7033), .I1(n7034), .O(\i16/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10994.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10995 (.I0(\rx_fifo/wr_index[1] ), .I1(\rx_fifo/wr_index[3] ), 
            .I2(\rx_fifo/wr_index[4] ), .I3(\rx_fifo/wr_index[2] ), .O(n7035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10995.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10996 (.I0(n7030), .I1(n7035), .O(\i16/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10996.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10997 (.I0(n7033), .I1(n7035), .O(\i16/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10997.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10998 (.I0(\rx_fifo/wr_index[3] ), .I1(\rx_fifo/wr_index[4] ), 
            .I2(\rx_fifo/wr_index[1] ), .I3(\rx_fifo/wr_index[2] ), .O(n7036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10998.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10999 (.I0(n7030), .I1(n7036), .O(\i16/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10999.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11000 (.I0(n7033), .I1(n7036), .O(\i16/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11000.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11001 (.I0(\rx_fifo/wr_index[1] ), .I1(\rx_fifo/wr_index[2] ), 
            .I2(\rx_fifo/wr_index[4] ), .I3(\rx_fifo/wr_index[3] ), .O(n7037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11001.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11002 (.I0(n7030), .I1(n7037), .O(\i16/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11002.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11003 (.I0(n7033), .I1(n7037), .O(\i16/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11003.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11004 (.I0(\rx_fifo/wr_index[2] ), .I1(\rx_fifo/wr_index[4] ), 
            .I2(\rx_fifo/wr_index[3] ), .I3(\rx_fifo/wr_index[1] ), .O(n7038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11004.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11005 (.I0(n7030), .I1(n7038), .O(\i16/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11005.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11006 (.I0(n7033), .I1(n7038), .O(\i16/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11006.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11007 (.I0(\rx_fifo/wr_index[1] ), .I1(\rx_fifo/wr_index[4] ), 
            .I2(\rx_fifo/wr_index[3] ), .I3(\rx_fifo/wr_index[2] ), .O(n7039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11007.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11008 (.I0(n7030), .I1(n7039), .O(\i16/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11008.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11009 (.I0(n7033), .I1(n7039), .O(\i16/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11009.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11010 (.I0(\rx_fifo/wr_index[4] ), .I1(\rx_fifo/wr_index[2] ), 
            .I2(\rx_fifo/wr_index[3] ), .I3(\rx_fifo/wr_index[1] ), .O(n7040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__11010.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__11011 (.I0(n7030), .I1(n7040), .O(\i16/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11011.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11012 (.I0(n7033), .I1(n7040), .O(\i16/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11012.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11013 (.I0(\rx_fifo/wr_index[1] ), .I1(\rx_fifo/wr_index[2] ), 
            .I2(\rx_fifo/wr_index[3] ), .I3(\rx_fifo/wr_index[4] ), .O(n7041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11013.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11014 (.I0(n7030), .I1(n7041), .O(\i16/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11014.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11015 (.I0(n7033), .I1(n7041), .O(\i16/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11015.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11016 (.I0(\rx_fifo/wr_index[2] ), .I1(\rx_fifo/wr_index[3] ), 
            .I2(\rx_fifo/wr_index[1] ), .I3(\rx_fifo/wr_index[4] ), .O(n7042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11016.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11017 (.I0(n7030), .I1(n7042), .O(\i16/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11017.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11018 (.I0(n7033), .I1(n7042), .O(\i16/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11018.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11019 (.I0(\rx_fifo/wr_index[1] ), .I1(\rx_fifo/wr_index[3] ), 
            .I2(\rx_fifo/wr_index[2] ), .I3(\rx_fifo/wr_index[4] ), .O(n7043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11019.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11020 (.I0(n7030), .I1(n7043), .O(\i16/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11020.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11021 (.I0(n7033), .I1(n7043), .O(\i16/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11021.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11022 (.I0(\rx_fifo/wr_index[3] ), .I1(\rx_fifo/wr_index[2] ), 
            .I2(\rx_fifo/wr_index[1] ), .I3(\rx_fifo/wr_index[4] ), .O(n7044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__11022.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__11023 (.I0(n7030), .I1(n7044), .O(\i16/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11023.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11024 (.I0(n7033), .I1(n7044), .O(\i16/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11024.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11025 (.I0(\rx_fifo/wr_index[1] ), .I1(\rx_fifo/wr_index[2] ), 
            .I2(\rx_fifo/wr_index[3] ), .I3(\rx_fifo/wr_index[4] ), .O(n7045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11025.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11026 (.I0(n7030), .I1(n7045), .O(\i16/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11026.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11027 (.I0(n7033), .I1(n7045), .O(\i16/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11027.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11028 (.I0(\rx_fifo/wr_index[2] ), .I1(\rx_fifo/wr_index[1] ), 
            .I2(\rx_fifo/wr_index[3] ), .I3(\rx_fifo/wr_index[4] ), .O(n7046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__11028.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__11029 (.I0(n7030), .I1(n7046), .O(\i16/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11029.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11030 (.I0(n7033), .I1(n7046), .O(\i16/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11030.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11031 (.I0(\rx_fifo/wr_index[1] ), .I1(\rx_fifo/wr_index[2] ), 
            .I2(\rx_fifo/wr_index[3] ), .I3(\rx_fifo/wr_index[4] ), .O(n7047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__11031.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__11032 (.I0(n7030), .I1(n7047), .O(\i16/n104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11032.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11033 (.I0(n7033), .I1(n7047), .O(\i16/n103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11033.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11034 (.I0(\rx_fifo/wr_index[1] ), .I1(\rx_fifo/wr_index[2] ), 
            .I2(\rx_fifo/wr_index[3] ), .I3(\rx_fifo/wr_index[4] ), .O(n7048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11034.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11035 (.I0(n7030), .I1(n7048), .O(\i16/n102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11035.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11036 (.I0(n7033), .I1(n7048), .O(\i16/n101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11036.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11037 (.I0(\rx_fifo/wr_index[6] ), .I1(\rx_fifo/wr_index[5] ), 
            .I2(n7029), .O(n7049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11037.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11038 (.I0(n7049), .I1(n7031), .O(\i16/n100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11038.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11039 (.I0(\rx_fifo/wr_index[6] ), .I1(\rx_fifo/wr_index[5] ), 
            .I2(n7032), .O(n7050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11039.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11040 (.I0(n7050), .I1(n7031), .O(\i16/n99 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11040.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11041 (.I0(n7049), .I1(n7034), .O(\i16/n98 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11041.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11042 (.I0(n7050), .I1(n7034), .O(\i16/n97 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11042.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11043 (.I0(n7049), .I1(n7035), .O(\i16/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11043.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11044 (.I0(n7050), .I1(n7035), .O(\i16/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11044.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11045 (.I0(n7049), .I1(n7036), .O(\i16/n94 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11045.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11046 (.I0(n7050), .I1(n7036), .O(\i16/n93 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11046.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11047 (.I0(n7049), .I1(n7037), .O(\i16/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11047.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11048 (.I0(n7050), .I1(n7037), .O(\i16/n91 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11048.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11049 (.I0(n7049), .I1(n7038), .O(\i16/n90 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11049.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11050 (.I0(n7050), .I1(n7038), .O(\i16/n89 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11050.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11051 (.I0(n7049), .I1(n7039), .O(\i16/n88 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11051.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11052 (.I0(n7050), .I1(n7039), .O(\i16/n87 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11052.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11053 (.I0(n7049), .I1(n7040), .O(\i16/n86 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11053.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11054 (.I0(n7050), .I1(n7040), .O(\i16/n85 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11054.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11055 (.I0(n7049), .I1(n7041), .O(\i16/n84 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11055.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11056 (.I0(n7050), .I1(n7041), .O(\i16/n83 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11056.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11057 (.I0(n7049), .I1(n7042), .O(\i16/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11057.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11058 (.I0(n7050), .I1(n7042), .O(\i16/n81 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11058.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11059 (.I0(n7049), .I1(n7043), .O(\i16/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11059.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11060 (.I0(n7050), .I1(n7043), .O(\i16/n79 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11060.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11061 (.I0(n7049), .I1(n7044), .O(\i16/n78 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11061.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11062 (.I0(n7050), .I1(n7044), .O(\i16/n77 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11062.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11063 (.I0(n7049), .I1(n7045), .O(\i16/n76 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11063.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11064 (.I0(n7050), .I1(n7045), .O(\i16/n75 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11064.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11065 (.I0(n7049), .I1(n7046), .O(\i16/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11065.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11066 (.I0(n7050), .I1(n7046), .O(\i16/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11066.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11067 (.I0(n7049), .I1(n7047), .O(\i16/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11067.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11068 (.I0(n7050), .I1(n7047), .O(\i16/n71 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11068.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11069 (.I0(n7049), .I1(n7048), .O(\i16/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11069.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11070 (.I0(n7050), .I1(n7048), .O(\i16/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11070.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11071 (.I0(\rx_fifo/wr_index[5] ), .I1(n7029), .I2(\rx_fifo/wr_index[6] ), 
            .O(n7051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11071.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11072 (.I0(n7051), .I1(n7031), .O(\i16/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11072.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11073 (.I0(\rx_fifo/wr_index[5] ), .I1(n7032), .I2(\rx_fifo/wr_index[6] ), 
            .O(n7052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11073.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11074 (.I0(n7052), .I1(n7031), .O(\i16/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11074.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11075 (.I0(n7051), .I1(n7034), .O(\i16/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11075.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11076 (.I0(n7052), .I1(n7034), .O(\i16/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11076.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11077 (.I0(n7051), .I1(n7035), .O(\i16/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11077.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11078 (.I0(n7052), .I1(n7035), .O(\i16/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11078.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11079 (.I0(n7051), .I1(n7036), .O(\i16/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11079.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11080 (.I0(n7052), .I1(n7036), .O(\i16/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11080.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11081 (.I0(n7051), .I1(n7037), .O(\i16/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11081.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11082 (.I0(n7052), .I1(n7037), .O(\i16/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11082.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11083 (.I0(n7051), .I1(n7038), .O(\i16/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11083.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11084 (.I0(n7052), .I1(n7038), .O(\i16/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11084.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11085 (.I0(n7051), .I1(n7039), .O(\i16/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11085.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11086 (.I0(n7052), .I1(n7039), .O(\i16/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11086.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11087 (.I0(n7051), .I1(n7040), .O(\i16/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11087.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11088 (.I0(n7052), .I1(n7040), .O(\i16/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11088.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11089 (.I0(n7051), .I1(n7041), .O(\i16/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11089.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11090 (.I0(n7052), .I1(n7041), .O(\i16/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11090.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11091 (.I0(n7051), .I1(n7042), .O(\i16/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11091.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11092 (.I0(n7052), .I1(n7042), .O(\i16/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11092.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11093 (.I0(n7051), .I1(n7043), .O(\i16/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11093.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11094 (.I0(n7052), .I1(n7043), .O(\i16/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11094.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11095 (.I0(n7051), .I1(n7044), .O(\i16/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11095.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11096 (.I0(n7052), .I1(n7044), .O(\i16/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11096.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11097 (.I0(n7051), .I1(n7045), .O(\i16/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11097.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11098 (.I0(n7052), .I1(n7045), .O(\i16/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11098.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11099 (.I0(n7051), .I1(n7046), .O(\i16/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11099.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11100 (.I0(n7052), .I1(n7046), .O(\i16/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11100.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11101 (.I0(n7051), .I1(n7047), .O(\i16/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11101.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11102 (.I0(n7052), .I1(n7047), .O(\i16/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11102.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11103 (.I0(n7051), .I1(n7048), .O(\i16/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11103.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11104 (.I0(n7052), .I1(n7048), .O(\i16/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11104.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11105 (.I0(n7029), .I1(\rx_fifo/wr_index[5] ), .I2(\rx_fifo/wr_index[6] ), 
            .O(n7053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11105.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11106 (.I0(n7053), .I1(n7031), .O(\i16/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11106.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11107 (.I0(n7032), .I1(\rx_fifo/wr_index[5] ), .I2(\rx_fifo/wr_index[6] ), 
            .O(n7054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11107.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11108 (.I0(n7054), .I1(n7031), .O(\i16/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11108.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11109 (.I0(n7053), .I1(n7034), .O(\i16/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11109.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11110 (.I0(n7054), .I1(n7034), .O(\i16/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11110.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11111 (.I0(n7053), .I1(n7035), .O(\i16/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11111.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11112 (.I0(n7054), .I1(n7035), .O(\i16/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11112.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11113 (.I0(n7053), .I1(n7036), .O(\i16/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11113.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11114 (.I0(n7054), .I1(n7036), .O(\i16/n29 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11114.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11115 (.I0(n7053), .I1(n7037), .O(\i16/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11115.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11116 (.I0(n7054), .I1(n7037), .O(\i16/n27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11116.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11117 (.I0(n7053), .I1(n7038), .O(\i16/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11117.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11118 (.I0(n7054), .I1(n7038), .O(\i16/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11118.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11119 (.I0(n7053), .I1(n7039), .O(\i16/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11119.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11120 (.I0(n7054), .I1(n7039), .O(\i16/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11120.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11121 (.I0(n7053), .I1(n7040), .O(\i16/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11121.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11122 (.I0(n7054), .I1(n7040), .O(\i16/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11122.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11123 (.I0(n7053), .I1(n7041), .O(\i16/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11123.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11124 (.I0(n7054), .I1(n7041), .O(\i16/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11124.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11125 (.I0(n7053), .I1(n7042), .O(\i16/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11125.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11126 (.I0(n7054), .I1(n7042), .O(\i16/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11126.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11127 (.I0(n7053), .I1(n7043), .O(\i16/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11127.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11128 (.I0(n7054), .I1(n7043), .O(\i16/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11128.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11129 (.I0(n7053), .I1(n7044), .O(\i16/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11129.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11130 (.I0(n7054), .I1(n7044), .O(\i16/n13 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11130.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11131 (.I0(n7053), .I1(n7045), .O(\i16/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11131.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11132 (.I0(n7054), .I1(n7045), .O(\i16/n11 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11132.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11133 (.I0(n7053), .I1(n7046), .O(\i16/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11133.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11134 (.I0(n7054), .I1(n7046), .O(\i16/n9 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11134.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11135 (.I0(n7053), .I1(n7047), .O(\i16/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11135.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11136 (.I0(n7054), .I1(n7047), .O(\i16/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11136.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11137 (.I0(n7053), .I1(n7048), .O(\i16/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11137.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11138 (.I0(n7054), .I1(n7048), .O(\i16/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11138.LUTMASK = 16'h8888;
    EFX_GBUFCE CLKBUF__1 (.CE(1'b1), .I(pll_clk), .O(\pll_clk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__1.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(tx_slowclk), .O(\tx_slowclk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__tx_dac_fsm_inst/add_18/i2  (.I0(\tx_dac_fsm_inst/sym_ctr[0] ), 
            .I1(1'b1), .CI(1'b0), .CO(n7059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(95)
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/add_18/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/add_18/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__tx_dac_fsm_inst/sub_20/add_2/i4  (.I0(\tx_dac_fsm_inst/sym_ctr[2] ), 
            .I1(1'b1), .CI(1'b0), .CO(n7058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(97)
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/sub_20/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/sub_20/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__tx_dac_fsm_inst/sub_20/add_2/i5  (.I0(n4167), .I1(1'b1), 
            .CI(1'b0), .CO(n7057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(97)
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/sub_20/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/sub_20/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__tx_dac_fsm_inst/add_129/i4  (.I0(n4161), .I1(1'b1), 
            .CI(1'b0), .CO(n7056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(197)
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/add_129/i4 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/add_129/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__tx_dac_fsm_inst/add_136/i4  (.I0(n4152), .I1(1'b1), 
            .CI(1'b0), .CO(n7055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Capstone\WES207\rtl\WES207_basic\rtl\tx_dac_fsm.sv(208)
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/add_136/i4 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__tx_dac_fsm_inst/add_136/i4 .I1_POLARITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_dfe71ff1_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_dfe71ff1_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_dfe71ff1_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_dfe71ff1_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_dfe71ff1_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_dfe71ff1_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_dfe71ff1_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_dfe71ff1_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_dfe71ff1_0
// module not written out since it is a black box. 
//

